-- from http://help.latticesemi.com/docs/webhelp/eng/wwhelp/wwhimpl/common/html/wwhelp.htm#href=Design%20Entry/inferring_ram_dual_port.htm
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
 
entity font_lb_dp_ram is
generic (
	addr_width : natural;
	data_width : natural);
port (
	addra_i	: in std_logic_vector (addr_width - 1 downto 0);
	wea_i	: in std_logic;
	clka_i	: in std_logic;
	dina_i	: in std_logic_vector (data_width - 1 downto 0);
	douta_o	: out std_logic_vector (data_width - 1 downto 0);
	addrb_i	: in std_logic_vector (addr_width - 1 downto 0);
	web_i	: in std_logic;
	clkb_i	: in std_logic;
	dinb_i	: in std_logic_vector (data_width - 1 downto 0);
	doutb_o	: out std_logic_vector (data_width - 1 downto 0));
end font_lb_dp_ram;
 
architecture rtl of font_lb_dp_ram is
	type mem_type is array ((2** addr_width) - 1 downto 0) of 
	std_logic_vector(data_width - 1 downto 0);
	signal mem : mem_type := (
-- odd lines (lower byte)
-- char 0x00='\0' 
--   =>	"00000000",	-- ........
   0 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
   1 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
   2 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
   3 =>	"00000000",	-- ........

-- char 0x01='\x01
--   =>	"01111110",	-- .######.
   4 =>	"10000001",	-- #......#
--   =>	"10100101",	-- #.#..#.#
   5 =>	"10000001",	-- #......#
--   =>	"10111101",	-- #.####.#
   6 =>	"10011001",	-- #..##..#
--   =>	"10000001",	-- #......#
   7 =>	"01111110",	-- .######.

-- char 0x02='\x02
--   =>	"01111110",	-- .######.
   8 =>	"11111111",	-- ########
--   =>	"11011011",	-- ##.##.##
   9 =>	"11111111",	-- ########
--   =>	"11000011",	-- ##....##
  10 =>	"11100111",	-- ###..###
--   =>	"11111111",	-- ########
  11 =>	"01111110",	-- .######.

-- char 0x03='\x03
--   =>	"01101100",	-- .##.##..
  12 =>	"11111110",	-- #######.
--   =>	"11111110",	-- #######.
  13 =>	"11111110",	-- #######.
--   =>	"01111100",	-- .#####..
  14 =>	"00111000",	-- ..###...
--   =>	"00010000",	-- ...#....
  15 =>	"00000000",	-- ........

-- char 0x04='\x04
--   =>	"00010000",	-- ...#....
  16 =>	"00111000",	-- ..###...
--   =>	"01111100",	-- .#####..
  17 =>	"11111110",	-- #######.
--   =>	"01111100",	-- .#####..
  18 =>	"00111000",	-- ..###...
--   =>	"00010000",	-- ...#....
  19 =>	"00000000",	-- ........

-- char 0x05='\x05
--   =>	"00111000",	-- ..###...
  20 =>	"01111100",	-- .#####..
--   =>	"00111000",	-- ..###...
  21 =>	"11111110",	-- #######.
--   =>	"11111110",	-- #######.
  22 =>	"11010110",	-- ##.#.##.
--   =>	"00010000",	-- ...#....
  23 =>	"00111000",	-- ..###...

-- char 0x06='\x06
--   =>	"00010000",	-- ...#....
  24 =>	"00010000",	-- ...#....
--   =>	"00111000",	-- ..###...
  25 =>	"01111100",	-- .#####..
--   =>	"11111110",	-- #######.
  26 =>	"01111100",	-- .#####..
--   =>	"00010000",	-- ...#....
  27 =>	"00111000",	-- ..###...

-- char 0x07='\a' 
--   =>	"00000000",	-- ........
  28 =>	"00000000",	-- ........
--   =>	"00011000",	-- ...##...
  29 =>	"00111100",	-- ..####..
--   =>	"00111100",	-- ..####..
  30 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........
  31 =>	"00000000",	-- ........

-- char 0x08='\b' 
--   =>	"11111111",	-- ########
  32 =>	"11111111",	-- ########
--   =>	"11100111",	-- ###..###
  33 =>	"11000011",	-- ##....##
--   =>	"11000011",	-- ##....##
  34 =>	"11100111",	-- ###..###
--   =>	"11111111",	-- ########
  35 =>	"11111111",	-- ########

-- char 0x09='\t' 
--   =>	"00000000",	-- ........
  36 =>	"00111100",	-- ..####..
--   =>	"01100110",	-- .##..##.
  37 =>	"01000010",	-- .#....#.
--   =>	"01000010",	-- .#....#.
  38 =>	"01100110",	-- .##..##.
--   =>	"00111100",	-- ..####..
  39 =>	"00000000",	-- ........

-- char 0x0a='\n' 
--   =>	"11111111",	-- ########
  40 =>	"11000011",	-- ##....##
--   =>	"10011001",	-- #..##..#
  41 =>	"10111101",	-- #.####.#
--   =>	"10111101",	-- #.####.#
  42 =>	"10011001",	-- #..##..#
--   =>	"11000011",	-- ##....##
  43 =>	"11111111",	-- ########

-- char 0x0b='\v' 
--   =>	"00001111",	-- ....####
  44 =>	"00000111",	-- .....###
--   =>	"00001111",	-- ....####
  45 =>	"01111101",	-- .#####.#
--   =>	"11001100",	-- ##..##..
  46 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
  47 =>	"01111000",	-- .####...

-- char 0x0c='\f' 
--   =>	"00111100",	-- ..####..
  48 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
  49 =>	"01100110",	-- .##..##.
--   =>	"00111100",	-- ..####..
  50 =>	"00011000",	-- ...##...
--   =>	"01111110",	-- .######.
  51 =>	"00011000",	-- ...##...

-- char 0x0d='\r' 
--   =>	"00111111",	-- ..######
  52 =>	"00110011",	-- ..##..##
--   =>	"00111111",	-- ..######
  53 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
  54 =>	"01110000",	-- .###....
--   =>	"11110000",	-- ####....
  55 =>	"11100000",	-- ###.....

-- char 0x0e='\x0e
--   =>	"01111111",	-- .#######
  56 =>	"01100011",	-- .##...##
--   =>	"01111111",	-- .#######
  57 =>	"01100011",	-- .##...##
--   =>	"01100011",	-- .##...##
  58 =>	"01100111",	-- .##..###
--   =>	"11100110",	-- ###..##.
  59 =>	"11000000",	-- ##......

-- char 0x0f='\x0f
--   =>	"00011000",	-- ...##...
  60 =>	"11011011",	-- ##.##.##
--   =>	"00111100",	-- ..####..
  61 =>	"11100111",	-- ###..###
--   =>	"11100111",	-- ###..###
  62 =>	"00111100",	-- ..####..
--   =>	"11011011",	-- ##.##.##
  63 =>	"00011000",	-- ...##...

-- char 0x10='\x10
--   =>	"10000000",	-- #.......
  64 =>	"11100000",	-- ###.....
--   =>	"11111000",	-- #####...
  65 =>	"11111110",	-- #######.
--   =>	"11111000",	-- #####...
  66 =>	"11100000",	-- ###.....
--   =>	"10000000",	-- #.......
  67 =>	"00000000",	-- ........

-- char 0x11='\x11
--   =>	"00000010",	-- ......#.
  68 =>	"00001110",	-- ....###.
--   =>	"00111110",	-- ..#####.
  69 =>	"11111110",	-- #######.
--   =>	"00111110",	-- ..#####.
  70 =>	"00001110",	-- ....###.
--   =>	"00000010",	-- ......#.
  71 =>	"00000000",	-- ........

-- char 0x12='\x12
--   =>	"00011000",	-- ...##...
  72 =>	"00111100",	-- ..####..
--   =>	"01111110",	-- .######.
  73 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
  74 =>	"01111110",	-- .######.
--   =>	"00111100",	-- ..####..
  75 =>	"00011000",	-- ...##...

-- char 0x13='\x13
--   =>	"01100110",	-- .##..##.
  76 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
  77 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
  78 =>	"00000000",	-- ........
--   =>	"01100110",	-- .##..##.
  79 =>	"00000000",	-- ........

-- char 0x14='\x14
--   =>	"01111111",	-- .#######
  80 =>	"11011011",	-- ##.##.##
--   =>	"11011011",	-- ##.##.##
  81 =>	"01111011",	-- .####.##
--   =>	"00011011",	-- ...##.##
  82 =>	"00011011",	-- ...##.##
--   =>	"00011011",	-- ...##.##
  83 =>	"00000000",	-- ........

-- char 0x15='\x15
--   =>	"00111110",	-- ..#####.
  84 =>	"01100011",	-- .##...##
--   =>	"00111000",	-- ..###...
  85 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
  86 =>	"00111000",	-- ..###...
--   =>	"11001100",	-- ##..##..
  87 =>	"01111000",	-- .####...

-- char 0x16='\x16
--   =>	"00000000",	-- ........
  88 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
  89 =>	"00000000",	-- ........
--   =>	"01111110",	-- .######.
  90 =>	"01111110",	-- .######.
--   =>	"01111110",	-- .######.
  91 =>	"00000000",	-- ........

-- char 0x17='\x17
--   =>	"00011000",	-- ...##...
  92 =>	"00111100",	-- ..####..
--   =>	"01111110",	-- .######.
  93 =>	"00011000",	-- ...##...
--   =>	"01111110",	-- .######.
  94 =>	"00111100",	-- ..####..
--   =>	"00011000",	-- ...##...
  95 =>	"11111111",	-- ########

-- char 0x18='\x18
--   =>	"00011000",	-- ...##...
  96 =>	"00111100",	-- ..####..
--   =>	"01111110",	-- .######.
  97 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
  98 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
  99 =>	"00000000",	-- ........

-- char 0x19='\x19
--   =>	"00011000",	-- ...##...
 100 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 101 =>	"00011000",	-- ...##...
--   =>	"01111110",	-- .######.
 102 =>	"00111100",	-- ..####..
--   =>	"00011000",	-- ...##...
 103 =>	"00000000",	-- ........

-- char 0x1a='\x1a
--   =>	"00000000",	-- ........
 104 =>	"00011000",	-- ...##...
--   =>	"00001100",	-- ....##..
 105 =>	"11111110",	-- #######.
--   =>	"00001100",	-- ....##..
 106 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........
 107 =>	"00000000",	-- ........

-- char 0x1b='\x1b
--   =>	"00000000",	-- ........
 108 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
 109 =>	"11111110",	-- #######.
--   =>	"01100000",	-- .##.....
 110 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 111 =>	"00000000",	-- ........

-- char 0x1c='\x1c
--   =>	"00000000",	-- ........
 112 =>	"00000000",	-- ........
--   =>	"11000000",	-- ##......
 113 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 114 =>	"11111110",	-- #######.
--   =>	"00000000",	-- ........
 115 =>	"00000000",	-- ........

-- char 0x1d='\x1d
--   =>	"00000000",	-- ........
 116 =>	"00100100",	-- ..#..#..
--   =>	"01100110",	-- .##..##.
 117 =>	"11111111",	-- ########
--   =>	"01100110",	-- .##..##.
 118 =>	"00100100",	-- ..#..#..
--   =>	"00000000",	-- ........
 119 =>	"00000000",	-- ........

-- char 0x1e='\x1e
--   =>	"00000000",	-- ........
 120 =>	"00011000",	-- ...##...
--   =>	"00111100",	-- ..####..
 121 =>	"01111110",	-- .######.
--   =>	"11111111",	-- ########
 122 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 123 =>	"00000000",	-- ........

-- char 0x1f='\x1f
--   =>	"00000000",	-- ........
 124 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 125 =>	"01111110",	-- .######.
--   =>	"00111100",	-- ..####..
 126 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........
 127 =>	"00000000",	-- ........

-- char 0x20=' '  
--   =>	"00000000",	-- ........
 128 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 129 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 130 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 131 =>	"00000000",	-- ........

-- char 0x21='!'  
--   =>	"00110000",	-- ..##....
 132 =>	"01111000",	-- .####...
--   =>	"01111000",	-- .####...
 133 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 134 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 135 =>	"00000000",	-- ........

-- char 0x22='\'' 
--   =>	"01101100",	-- .##.##..
 136 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 137 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 138 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 139 =>	"00000000",	-- ........

-- char 0x23='#'  
--   =>	"01101100",	-- .##.##..
 140 =>	"01101100",	-- .##.##..
--   =>	"11111110",	-- #######.
 141 =>	"01101100",	-- .##.##..
--   =>	"11111110",	-- #######.
 142 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 143 =>	"00000000",	-- ........

-- char 0x24='$'  
--   =>	"00110000",	-- ..##....
 144 =>	"01111100",	-- .#####..
--   =>	"11000000",	-- ##......
 145 =>	"01111000",	-- .####...
--   =>	"00001100",	-- ....##..
 146 =>	"11111000",	-- #####...
--   =>	"00110000",	-- ..##....
 147 =>	"00000000",	-- ........

-- char 0x25='%'  
--   =>	"00000000",	-- ........
 148 =>	"11000110",	-- ##...##.
--   =>	"11001100",	-- ##..##..
 149 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
 150 =>	"01100110",	-- .##..##.
--   =>	"11000110",	-- ##...##.
 151 =>	"00000000",	-- ........

-- char 0x26='&'  
--   =>	"00111000",	-- ..###...
 152 =>	"01101100",	-- .##.##..
--   =>	"00111000",	-- ..###...
 153 =>	"01110110",	-- .###.##.
--   =>	"11011100",	-- ##.###..
 154 =>	"11001100",	-- ##..##..
--   =>	"01110110",	-- .###.##.
 155 =>	"00000000",	-- ........

-- char 0x27='\"' 
--   =>	"01100000",	-- .##.....
 156 =>	"01100000",	-- .##.....
--   =>	"11000000",	-- ##......
 157 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 158 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 159 =>	"00000000",	-- ........

-- char 0x28='('  
--   =>	"00011000",	-- ...##...
 160 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
 161 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 162 =>	"00110000",	-- ..##....
--   =>	"00011000",	-- ...##...
 163 =>	"00000000",	-- ........

-- char 0x29=')'  
--   =>	"01100000",	-- .##.....
 164 =>	"00110000",	-- ..##....
--   =>	"00011000",	-- ...##...
 165 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 166 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
 167 =>	"00000000",	-- ........

-- char 0x2a='*'  
--   =>	"00000000",	-- ........
 168 =>	"01100110",	-- .##..##.
--   =>	"00111100",	-- ..####..
 169 =>	"11111111",	-- ########
--   =>	"00111100",	-- ..####..
 170 =>	"01100110",	-- .##..##.
--   =>	"00000000",	-- ........
 171 =>	"00000000",	-- ........

-- char 0x2b='+'  
--   =>	"00000000",	-- ........
 172 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 173 =>	"11111100",	-- ######..
--   =>	"00110000",	-- ..##....
 174 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 175 =>	"00000000",	-- ........

-- char 0x2c=','  
--   =>	"00000000",	-- ........
 176 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 177 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 178 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 179 =>	"01100000",	-- .##.....

-- char 0x2d='-'  
--   =>	"00000000",	-- ........
 180 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 181 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........
 182 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 183 =>	"00000000",	-- ........

-- char 0x2e='.'  
--   =>	"00000000",	-- ........
 184 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 185 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 186 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 187 =>	"00000000",	-- ........

-- char 0x2f='/'  
--   =>	"00000110",	-- .....##.
 188 =>	"00001100",	-- ....##..
--   =>	"00011000",	-- ...##...
 189 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
 190 =>	"11000000",	-- ##......
--   =>	"10000000",	-- #.......
 191 =>	"00000000",	-- ........

-- char 0x30='0'  
--   =>	"01111100",	-- .#####..
 192 =>	"11000110",	-- ##...##.
--   =>	"11001110",	-- ##..###.
 193 =>	"11011110",	-- ##.####.
--   =>	"11110110",	-- ####.##.
 194 =>	"11100110",	-- ###..##.
--   =>	"01111100",	-- .#####..
 195 =>	"00000000",	-- ........

-- char 0x31='1'  
--   =>	"00110000",	-- ..##....
 196 =>	"01110000",	-- .###....
--   =>	"00110000",	-- ..##....
 197 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 198 =>	"00110000",	-- ..##....
--   =>	"11111100",	-- ######..
 199 =>	"00000000",	-- ........

-- char 0x32='2'  
--   =>	"01111000",	-- .####...
 200 =>	"11001100",	-- ##..##..
--   =>	"00001100",	-- ....##..
 201 =>	"00111000",	-- ..###...
--   =>	"01100000",	-- .##.....
 202 =>	"11001100",	-- ##..##..
--   =>	"11111100",	-- ######..
 203 =>	"00000000",	-- ........

-- char 0x33='3'  
--   =>	"01111000",	-- .####...
 204 =>	"11001100",	-- ##..##..
--   =>	"00001100",	-- ....##..
 205 =>	"00111000",	-- ..###...
--   =>	"00001100",	-- ....##..
 206 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 207 =>	"00000000",	-- ........

-- char 0x34='4'  
--   =>	"00011100",	-- ...###..
 208 =>	"00111100",	-- ..####..
--   =>	"01101100",	-- .##.##..
 209 =>	"11001100",	-- ##..##..
--   =>	"11111110",	-- #######.
 210 =>	"00001100",	-- ....##..
--   =>	"00011110",	-- ...####.
 211 =>	"00000000",	-- ........

-- char 0x35='5'  
--   =>	"11111100",	-- ######..
 212 =>	"11000000",	-- ##......
--   =>	"11111000",	-- #####...
 213 =>	"00001100",	-- ....##..
--   =>	"00001100",	-- ....##..
 214 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 215 =>	"00000000",	-- ........

-- char 0x36='6'  
--   =>	"00111000",	-- ..###...
 216 =>	"01100000",	-- .##.....
--   =>	"11000000",	-- ##......
 217 =>	"11111000",	-- #####...
--   =>	"11001100",	-- ##..##..
 218 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 219 =>	"00000000",	-- ........

-- char 0x37='7'  
--   =>	"11111100",	-- ######..
 220 =>	"11001100",	-- ##..##..
--   =>	"00001100",	-- ....##..
 221 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
 222 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 223 =>	"00000000",	-- ........

-- char 0x38='8'  
--   =>	"01111000",	-- .####...
 224 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 225 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 226 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 227 =>	"00000000",	-- ........

-- char 0x39='9'  
--   =>	"01111000",	-- .####...
 228 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 229 =>	"01111100",	-- .#####..
--   =>	"00001100",	-- ....##..
 230 =>	"00011000",	-- ...##...
--   =>	"01110000",	-- .###....
 231 =>	"00000000",	-- ........

-- char 0x3a=':'  
--   =>	"00000000",	-- ........
 232 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 233 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 234 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 235 =>	"00000000",	-- ........

-- char 0x3b=';'  
--   =>	"00000000",	-- ........
 236 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 237 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 238 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 239 =>	"01100000",	-- .##.....

-- char 0x3c='<'  
--   =>	"00011000",	-- ...##...
 240 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
 241 =>	"11000000",	-- ##......
--   =>	"01100000",	-- .##.....
 242 =>	"00110000",	-- ..##....
--   =>	"00011000",	-- ...##...
 243 =>	"00000000",	-- ........

-- char 0x3d='='  
--   =>	"00000000",	-- ........
 244 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 245 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 246 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........
 247 =>	"00000000",	-- ........

-- char 0x3e='>'  
--   =>	"01100000",	-- .##.....
 248 =>	"00110000",	-- ..##....
--   =>	"00011000",	-- ...##...
 249 =>	"00001100",	-- ....##..
--   =>	"00011000",	-- ...##...
 250 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
 251 =>	"00000000",	-- ........

-- char 0x3f='?'  
--   =>	"01111000",	-- .####...
 252 =>	"11001100",	-- ##..##..
--   =>	"00001100",	-- ....##..
 253 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
 254 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 255 =>	"00000000",	-- ........

-- char 0x40='@'  
--   =>	"01111100",	-- .#####..
 256 =>	"11000110",	-- ##...##.
--   =>	"11011110",	-- ##.####.
 257 =>	"11011110",	-- ##.####.
--   =>	"11011110",	-- ##.####.
 258 =>	"11000000",	-- ##......
--   =>	"01111000",	-- .####...
 259 =>	"00000000",	-- ........

-- char 0x41='A'  
--   =>	"00110000",	-- ..##....
 260 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 261 =>	"11001100",	-- ##..##..
--   =>	"11111100",	-- ######..
 262 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 263 =>	"00000000",	-- ........

-- char 0x42='B'  
--   =>	"11111100",	-- ######..
 264 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 265 =>	"01111100",	-- .#####..
--   =>	"01100110",	-- .##..##.
 266 =>	"01100110",	-- .##..##.
--   =>	"11111100",	-- ######..
 267 =>	"00000000",	-- ........

-- char 0x43='C'  
--   =>	"00111100",	-- ..####..
 268 =>	"01100110",	-- .##..##.
--   =>	"11000000",	-- ##......
 269 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 270 =>	"01100110",	-- .##..##.
--   =>	"00111100",	-- ..####..
 271 =>	"00000000",	-- ........

-- char 0x44='D'  
--   =>	"11111000",	-- #####...
 272 =>	"01101100",	-- .##.##..
--   =>	"01100110",	-- .##..##.
 273 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 274 =>	"01101100",	-- .##.##..
--   =>	"11111000",	-- #####...
 275 =>	"00000000",	-- ........

-- char 0x45='E'  
--   =>	"11111110",	-- #######.
 276 =>	"01100010",	-- .##...#.
--   =>	"01101000",	-- .##.#...
 277 =>	"01111000",	-- .####...
--   =>	"01101000",	-- .##.#...
 278 =>	"01100010",	-- .##...#.
--   =>	"11111110",	-- #######.
 279 =>	"00000000",	-- ........

-- char 0x46='F'  
--   =>	"11111110",	-- #######.
 280 =>	"01100010",	-- .##...#.
--   =>	"01101000",	-- .##.#...
 281 =>	"01111000",	-- .####...
--   =>	"01101000",	-- .##.#...
 282 =>	"01100000",	-- .##.....
--   =>	"11110000",	-- ####....
 283 =>	"00000000",	-- ........

-- char 0x47='G'  
--   =>	"00111100",	-- ..####..
 284 =>	"01100110",	-- .##..##.
--   =>	"11000000",	-- ##......
 285 =>	"11000000",	-- ##......
--   =>	"11001110",	-- ##..###.
 286 =>	"01100110",	-- .##..##.
--   =>	"00111110",	-- ..#####.
 287 =>	"00000000",	-- ........

-- char 0x48='H'  
--   =>	"11001100",	-- ##..##..
 288 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 289 =>	"11111100",	-- ######..
--   =>	"11001100",	-- ##..##..
 290 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 291 =>	"00000000",	-- ........

-- char 0x49='I'  
--   =>	"01111000",	-- .####...
 292 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 293 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 294 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 295 =>	"00000000",	-- ........

-- char 0x4a='J'  
--   =>	"00011110",	-- ...####.
 296 =>	"00001100",	-- ....##..
--   =>	"00001100",	-- ....##..
 297 =>	"00001100",	-- ....##..
--   =>	"11001100",	-- ##..##..
 298 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 299 =>	"00000000",	-- ........

-- char 0x4b='K'  
--   =>	"11100110",	-- ###..##.
 300 =>	"01100110",	-- .##..##.
--   =>	"01101100",	-- .##.##..
 301 =>	"01111000",	-- .####...
--   =>	"01101100",	-- .##.##..
 302 =>	"01100110",	-- .##..##.
--   =>	"11100110",	-- ###..##.
 303 =>	"00000000",	-- ........

-- char 0x4c='L'  
--   =>	"11110000",	-- ####....
 304 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 305 =>	"01100000",	-- .##.....
--   =>	"01100010",	-- .##...#.
 306 =>	"01100110",	-- .##..##.
--   =>	"11111110",	-- #######.
 307 =>	"00000000",	-- ........

-- char 0x4d='M'  
--   =>	"11000110",	-- ##...##.
 308 =>	"11101110",	-- ###.###.
--   =>	"11111110",	-- #######.
 309 =>	"11111110",	-- #######.
--   =>	"11010110",	-- ##.#.##.
 310 =>	"11000110",	-- ##...##.
--   =>	"11000110",	-- ##...##.
 311 =>	"00000000",	-- ........

-- char 0x4e='N'  
--   =>	"11000110",	-- ##...##.
 312 =>	"11100110",	-- ###..##.
--   =>	"11110110",	-- ####.##.
 313 =>	"11011110",	-- ##.####.
--   =>	"11001110",	-- ##..###.
 314 =>	"11000110",	-- ##...##.
--   =>	"11000110",	-- ##...##.
 315 =>	"00000000",	-- ........

-- char 0x4f='O'  
--   =>	"00111000",	-- ..###...
 316 =>	"01101100",	-- .##.##..
--   =>	"11000110",	-- ##...##.
 317 =>	"11000110",	-- ##...##.
--   =>	"11000110",	-- ##...##.
 318 =>	"01101100",	-- .##.##..
--   =>	"00111000",	-- ..###...
 319 =>	"00000000",	-- ........

-- char 0x50='P'  
--   =>	"11111100",	-- ######..
 320 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 321 =>	"01111100",	-- .#####..
--   =>	"01100000",	-- .##.....
 322 =>	"01100000",	-- .##.....
--   =>	"11110000",	-- ####....
 323 =>	"00000000",	-- ........

-- char 0x51='Q'  
--   =>	"01111000",	-- .####...
 324 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 325 =>	"11001100",	-- ##..##..
--   =>	"11011100",	-- ##.###..
 326 =>	"01111000",	-- .####...
--   =>	"00011100",	-- ...###..
 327 =>	"00000000",	-- ........

-- char 0x52='R'  
--   =>	"11111100",	-- ######..
 328 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 329 =>	"01111100",	-- .#####..
--   =>	"01101100",	-- .##.##..
 330 =>	"01100110",	-- .##..##.
--   =>	"11100110",	-- ###..##.
 331 =>	"00000000",	-- ........

-- char 0x53='S'  
--   =>	"01111000",	-- .####...
 332 =>	"11001100",	-- ##..##..
--   =>	"01100000",	-- .##.....
 333 =>	"00110000",	-- ..##....
--   =>	"00011000",	-- ...##...
 334 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 335 =>	"00000000",	-- ........

-- char 0x54='T'  
--   =>	"11111100",	-- ######..
 336 =>	"10110100",	-- #.##.#..
--   =>	"00110000",	-- ..##....
 337 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 338 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 339 =>	"00000000",	-- ........

-- char 0x55='U'  
--   =>	"11001100",	-- ##..##..
 340 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 341 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 342 =>	"11001100",	-- ##..##..
--   =>	"11111100",	-- ######..
 343 =>	"00000000",	-- ........

-- char 0x56='V'  
--   =>	"11001100",	-- ##..##..
 344 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 345 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 346 =>	"01111000",	-- .####...
--   =>	"00110000",	-- ..##....
 347 =>	"00000000",	-- ........

-- char 0x57='W'  
--   =>	"11000110",	-- ##...##.
 348 =>	"11000110",	-- ##...##.
--   =>	"11000110",	-- ##...##.
 349 =>	"11010110",	-- ##.#.##.
--   =>	"11111110",	-- #######.
 350 =>	"11101110",	-- ###.###.
--   =>	"11000110",	-- ##...##.
 351 =>	"00000000",	-- ........

-- char 0x58='X'  
--   =>	"11000110",	-- ##...##.
 352 =>	"11000110",	-- ##...##.
--   =>	"01101100",	-- .##.##..
 353 =>	"00111000",	-- ..###...
--   =>	"00111000",	-- ..###...
 354 =>	"01101100",	-- .##.##..
--   =>	"11000110",	-- ##...##.
 355 =>	"00000000",	-- ........

-- char 0x59='Y'  
--   =>	"11001100",	-- ##..##..
 356 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 357 =>	"01111000",	-- .####...
--   =>	"00110000",	-- ..##....
 358 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 359 =>	"00000000",	-- ........

-- char 0x5a='Z'  
--   =>	"11111110",	-- #######.
 360 =>	"11000110",	-- ##...##.
--   =>	"10001100",	-- #...##..
 361 =>	"00011000",	-- ...##...
--   =>	"00110010",	-- ..##..#.
 362 =>	"01100110",	-- .##..##.
--   =>	"11111110",	-- #######.
 363 =>	"00000000",	-- ........

-- char 0x5b='['  
--   =>	"01111000",	-- .####...
 364 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 365 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 366 =>	"01100000",	-- .##.....
--   =>	"01111000",	-- .####...
 367 =>	"00000000",	-- ........

-- char 0x5c='\\' 
--   =>	"11000000",	-- ##......
 368 =>	"01100000",	-- .##.....
--   =>	"00110000",	-- ..##....
 369 =>	"00011000",	-- ...##...
--   =>	"00001100",	-- ....##..
 370 =>	"00000110",	-- .....##.
--   =>	"00000010",	-- ......#.
 371 =>	"00000000",	-- ........

-- char 0x5d=']'  
--   =>	"01111000",	-- .####...
 372 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 373 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 374 =>	"00011000",	-- ...##...
--   =>	"01111000",	-- .####...
 375 =>	"00000000",	-- ........

-- char 0x5e='^'  
--   =>	"00010000",	-- ...#....
 376 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 377 =>	"11000110",	-- ##...##.
--   =>	"00000000",	-- ........
 378 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 379 =>	"00000000",	-- ........

-- char 0x5f='_'  
--   =>	"00000000",	-- ........
 380 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 381 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 382 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 383 =>	"11111111",	-- ########

-- char 0x60='`'  
--   =>	"00110000",	-- ..##....
 384 =>	"00110000",	-- ..##....
--   =>	"00011000",	-- ...##...
 385 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 386 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 387 =>	"00000000",	-- ........

-- char 0x61='a'  
--   =>	"00000000",	-- ........
 388 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 389 =>	"00001100",	-- ....##..
--   =>	"01111100",	-- .#####..
 390 =>	"11001100",	-- ##..##..
--   =>	"01110110",	-- .###.##.
 391 =>	"00000000",	-- ........

-- char 0x62='b'  
--   =>	"11100000",	-- ###.....
 392 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 393 =>	"01111100",	-- .#####..
--   =>	"01100110",	-- .##..##.
 394 =>	"01100110",	-- .##..##.
--   =>	"11011100",	-- ##.###..
 395 =>	"00000000",	-- ........

-- char 0x63='c'  
--   =>	"00000000",	-- ........
 396 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 397 =>	"11001100",	-- ##..##..
--   =>	"11000000",	-- ##......
 398 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 399 =>	"00000000",	-- ........

-- char 0x64='d'  
--   =>	"00011100",	-- ...###..
 400 =>	"00001100",	-- ....##..
--   =>	"00001100",	-- ....##..
 401 =>	"01111100",	-- .#####..
--   =>	"11001100",	-- ##..##..
 402 =>	"11001100",	-- ##..##..
--   =>	"01110110",	-- .###.##.
 403 =>	"00000000",	-- ........

-- char 0x65='e'  
--   =>	"00000000",	-- ........
 404 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 405 =>	"11001100",	-- ##..##..
--   =>	"11111100",	-- ######..
 406 =>	"11000000",	-- ##......
--   =>	"01111000",	-- .####...
 407 =>	"00000000",	-- ........

-- char 0x66='f'  
--   =>	"00111000",	-- ..###...
 408 =>	"01101100",	-- .##.##..
--   =>	"01100000",	-- .##.....
 409 =>	"11110000",	-- ####....
--   =>	"01100000",	-- .##.....
 410 =>	"01100000",	-- .##.....
--   =>	"11110000",	-- ####....
 411 =>	"00000000",	-- ........

-- char 0x67='g'  
--   =>	"00000000",	-- ........
 412 =>	"00000000",	-- ........
--   =>	"01110110",	-- .###.##.
 413 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 414 =>	"01111100",	-- .#####..
--   =>	"00001100",	-- ....##..
 415 =>	"11111000",	-- #####...

-- char 0x68='h'  
--   =>	"11100000",	-- ###.....
 416 =>	"01100000",	-- .##.....
--   =>	"01101100",	-- .##.##..
 417 =>	"01110110",	-- .###.##.
--   =>	"01100110",	-- .##..##.
 418 =>	"01100110",	-- .##..##.
--   =>	"11100110",	-- ###..##.
 419 =>	"00000000",	-- ........

-- char 0x69='i'  
--   =>	"00110000",	-- ..##....
 420 =>	"00000000",	-- ........
--   =>	"01110000",	-- .###....
 421 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 422 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 423 =>	"00000000",	-- ........

-- char 0x6a='j'  
--   =>	"00001100",	-- ....##..
 424 =>	"00000000",	-- ........
--   =>	"00001100",	-- ....##..
 425 =>	"00001100",	-- ....##..
--   =>	"00001100",	-- ....##..
 426 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 427 =>	"01111000",	-- .####...

-- char 0x6b='k'  
--   =>	"11100000",	-- ###.....
 428 =>	"01100000",	-- .##.....
--   =>	"01100110",	-- .##..##.
 429 =>	"01101100",	-- .##.##..
--   =>	"01111000",	-- .####...
 430 =>	"01101100",	-- .##.##..
--   =>	"11100110",	-- ###..##.
 431 =>	"00000000",	-- ........

-- char 0x6c='l'  
--   =>	"01110000",	-- .###....
 432 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 433 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 434 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 435 =>	"00000000",	-- ........

-- char 0x6d='m'  
--   =>	"00000000",	-- ........
 436 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 437 =>	"11111110",	-- #######.
--   =>	"11111110",	-- #######.
 438 =>	"11010110",	-- ##.#.##.
--   =>	"11000110",	-- ##...##.
 439 =>	"00000000",	-- ........

-- char 0x6e='n'  
--   =>	"00000000",	-- ........
 440 =>	"00000000",	-- ........
--   =>	"11111000",	-- #####...
 441 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 442 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 443 =>	"00000000",	-- ........

-- char 0x6f='o'  
--   =>	"00000000",	-- ........
 444 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 445 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 446 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 447 =>	"00000000",	-- ........

-- char 0x70='p'  
--   =>	"00000000",	-- ........
 448 =>	"00000000",	-- ........
--   =>	"11011100",	-- ##.###..
 449 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 450 =>	"01111100",	-- .#####..
--   =>	"01100000",	-- .##.....
 451 =>	"11110000",	-- ####....

-- char 0x71='q'  
--   =>	"00000000",	-- ........
 452 =>	"00000000",	-- ........
--   =>	"01110110",	-- .###.##.
 453 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 454 =>	"01111100",	-- .#####..
--   =>	"00001100",	-- ....##..
 455 =>	"00011110",	-- ...####.

-- char 0x72='r'  
--   =>	"00000000",	-- ........
 456 =>	"00000000",	-- ........
--   =>	"11011100",	-- ##.###..
 457 =>	"01110110",	-- .###.##.
--   =>	"01100110",	-- .##..##.
 458 =>	"01100000",	-- .##.....
--   =>	"11110000",	-- ####....
 459 =>	"00000000",	-- ........

-- char 0x73='s'  
--   =>	"00000000",	-- ........
 460 =>	"00000000",	-- ........
--   =>	"01111100",	-- .#####..
 461 =>	"11000000",	-- ##......
--   =>	"01111000",	-- .####...
 462 =>	"00001100",	-- ....##..
--   =>	"11111000",	-- #####...
 463 =>	"00000000",	-- ........

-- char 0x74='t'  
--   =>	"00010000",	-- ...#....
 464 =>	"00110000",	-- ..##....
--   =>	"01111100",	-- .#####..
 465 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 466 =>	"00110100",	-- ..##.#..
--   =>	"00011000",	-- ...##...
 467 =>	"00000000",	-- ........

-- char 0x75='u'  
--   =>	"00000000",	-- ........
 468 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 469 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 470 =>	"11001100",	-- ##..##..
--   =>	"01110110",	-- .###.##.
 471 =>	"00000000",	-- ........

-- char 0x76='v'  
--   =>	"00000000",	-- ........
 472 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 473 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 474 =>	"01111000",	-- .####...
--   =>	"00110000",	-- ..##....
 475 =>	"00000000",	-- ........

-- char 0x77='w'  
--   =>	"00000000",	-- ........
 476 =>	"00000000",	-- ........
--   =>	"11000110",	-- ##...##.
 477 =>	"11010110",	-- ##.#.##.
--   =>	"11111110",	-- #######.
 478 =>	"11111110",	-- #######.
--   =>	"01101100",	-- .##.##..
 479 =>	"00000000",	-- ........

-- char 0x78='x'  
--   =>	"00000000",	-- ........
 480 =>	"00000000",	-- ........
--   =>	"11000110",	-- ##...##.
 481 =>	"01101100",	-- .##.##..
--   =>	"00111000",	-- ..###...
 482 =>	"01101100",	-- .##.##..
--   =>	"11000110",	-- ##...##.
 483 =>	"00000000",	-- ........

-- char 0x79='y'  
--   =>	"00000000",	-- ........
 484 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 485 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 486 =>	"01111100",	-- .#####..
--   =>	"00001100",	-- ....##..
 487 =>	"11111000",	-- #####...

-- char 0x7a='z'  
--   =>	"00000000",	-- ........
 488 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 489 =>	"10011000",	-- #..##...
--   =>	"00110000",	-- ..##....
 490 =>	"01100100",	-- .##..#..
--   =>	"11111100",	-- ######..
 491 =>	"00000000",	-- ........

-- char 0x7b='{'  
--   =>	"00011100",	-- ...###..
 492 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 493 =>	"11100000",	-- ###.....
--   =>	"00110000",	-- ..##....
 494 =>	"00110000",	-- ..##....
--   =>	"00011100",	-- ...###..
 495 =>	"00000000",	-- ........

-- char 0x7c='|'  
--   =>	"00011000",	-- ...##...
 496 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 497 =>	"00000000",	-- ........
--   =>	"00011000",	-- ...##...
 498 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 499 =>	"00000000",	-- ........

-- char 0x7d='}'  
--   =>	"11100000",	-- ###.....
 500 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 501 =>	"00011100",	-- ...###..
--   =>	"00110000",	-- ..##....
 502 =>	"00110000",	-- ..##....
--   =>	"11100000",	-- ###.....
 503 =>	"00000000",	-- ........

-- char 0x7e='~'  
--   =>	"01110110",	-- .###.##.
 504 =>	"11011100",	-- ##.###..
--   =>	"00000000",	-- ........
 505 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 506 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 507 =>	"00000000",	-- ........

-- char 0x7f='\x7f
--   =>	"00000000",	-- ........
 508 =>	"00010000",	-- ...#....
--   =>	"00111000",	-- ..###...
 509 =>	"01101100",	-- .##.##..
--   =>	"11000110",	-- ##...##.
 510 =>	"11000110",	-- ##...##.
--   =>	"11111110",	-- #######.
 511 =>	"00000000",	-- ........

-- char 0x80='\x80
--   =>	"01111000",	-- .####...
 512 =>	"11001100",	-- ##..##..
--   =>	"11000000",	-- ##......
 513 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 514 =>	"00011000",	-- ...##...
--   =>	"00001100",	-- ....##..
 515 =>	"01111000",	-- .####...

-- char 0x81='\x81
--   =>	"00000000",	-- ........
 516 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........
 517 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 518 =>	"11001100",	-- ##..##..
--   =>	"01111110",	-- .######.
 519 =>	"00000000",	-- ........

-- char 0x82='\x82
--   =>	"00011100",	-- ...###..
 520 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 521 =>	"11001100",	-- ##..##..
--   =>	"11111100",	-- ######..
 522 =>	"11000000",	-- ##......
--   =>	"01111000",	-- .####...
 523 =>	"00000000",	-- ........

-- char 0x83='\x83
--   =>	"01111110",	-- .######.
 524 =>	"11000011",	-- ##....##
--   =>	"00111100",	-- ..####..
 525 =>	"00000110",	-- .....##.
--   =>	"00111110",	-- ..#####.
 526 =>	"01100110",	-- .##..##.
--   =>	"00111111",	-- ..######
 527 =>	"00000000",	-- ........

-- char 0x84='\x84
--   =>	"11001100",	-- ##..##..
 528 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 529 =>	"00001100",	-- ....##..
--   =>	"01111100",	-- .#####..
 530 =>	"11001100",	-- ##..##..
--   =>	"01111110",	-- .######.
 531 =>	"00000000",	-- ........

-- char 0x85='\x85
--   =>	"11100000",	-- ###.....
 532 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 533 =>	"00001100",	-- ....##..
--   =>	"01111100",	-- .#####..
 534 =>	"11001100",	-- ##..##..
--   =>	"01111110",	-- .######.
 535 =>	"00000000",	-- ........

-- char 0x86='\x86
--   =>	"00110000",	-- ..##....
 536 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 537 =>	"00001100",	-- ....##..
--   =>	"01111100",	-- .#####..
 538 =>	"11001100",	-- ##..##..
--   =>	"01111110",	-- .######.
 539 =>	"00000000",	-- ........

-- char 0x87='\x87
--   =>	"00000000",	-- ........
 540 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 541 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 542 =>	"01111000",	-- .####...
--   =>	"00001100",	-- ....##..
 543 =>	"00111000",	-- ..###...

-- char 0x88='\x88
--   =>	"01111110",	-- .######.
 544 =>	"11000011",	-- ##....##
--   =>	"00111100",	-- ..####..
 545 =>	"01100110",	-- .##..##.
--   =>	"01111110",	-- .######.
 546 =>	"01100000",	-- .##.....
--   =>	"00111100",	-- ..####..
 547 =>	"00000000",	-- ........

-- char 0x89='\x89
--   =>	"11001100",	-- ##..##..
 548 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 549 =>	"11001100",	-- ##..##..
--   =>	"11111100",	-- ######..
 550 =>	"11000000",	-- ##......
--   =>	"01111000",	-- .####...
 551 =>	"00000000",	-- ........

-- char 0x8a='\x8a
--   =>	"11100000",	-- ###.....
 552 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 553 =>	"11001100",	-- ##..##..
--   =>	"11111100",	-- ######..
 554 =>	"11000000",	-- ##......
--   =>	"01111000",	-- .####...
 555 =>	"00000000",	-- ........

-- char 0x8b='\x8b
--   =>	"11001100",	-- ##..##..
 556 =>	"00000000",	-- ........
--   =>	"01110000",	-- .###....
 557 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 558 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 559 =>	"00000000",	-- ........

-- char 0x8c='\x8c
--   =>	"01111100",	-- .#####..
 560 =>	"11000110",	-- ##...##.
--   =>	"00111000",	-- ..###...
 561 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 562 =>	"00011000",	-- ...##...
--   =>	"00111100",	-- ..####..
 563 =>	"00000000",	-- ........

-- char 0x8d='\x8d
--   =>	"11100000",	-- ###.....
 564 =>	"00000000",	-- ........
--   =>	"01110000",	-- .###....
 565 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 566 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 567 =>	"00000000",	-- ........

-- char 0x8e='\x8e
--   =>	"11000110",	-- ##...##.
 568 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 569 =>	"11000110",	-- ##...##.
--   =>	"11111110",	-- #######.
 570 =>	"11000110",	-- ##...##.
--   =>	"11000110",	-- ##...##.
 571 =>	"00000000",	-- ........

-- char 0x8f='\x8f
--   =>	"00110000",	-- ..##....
 572 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 573 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 574 =>	"11111100",	-- ######..
--   =>	"11001100",	-- ##..##..
 575 =>	"00000000",	-- ........

-- char 0x90='\x90
--   =>	"00011100",	-- ...###..
 576 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 577 =>	"01100000",	-- .##.....
--   =>	"01111000",	-- .####...
 578 =>	"01100000",	-- .##.....
--   =>	"11111100",	-- ######..
 579 =>	"00000000",	-- ........

-- char 0x91='\x91
--   =>	"00000000",	-- ........
 580 =>	"00000000",	-- ........
--   =>	"01111111",	-- .#######
 581 =>	"00001100",	-- ....##..
--   =>	"01111111",	-- .#######
 582 =>	"11001100",	-- ##..##..
--   =>	"01111111",	-- .#######
 583 =>	"00000000",	-- ........

-- char 0x92='\x92
--   =>	"00111110",	-- ..#####.
 584 =>	"01101100",	-- .##.##..
--   =>	"11001100",	-- ##..##..
 585 =>	"11111110",	-- #######.
--   =>	"11001100",	-- ##..##..
 586 =>	"11001100",	-- ##..##..
--   =>	"11001110",	-- ##..###.
 587 =>	"00000000",	-- ........

-- char 0x93='\x93
--   =>	"01111000",	-- .####...
 588 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........
 589 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 590 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 591 =>	"00000000",	-- ........

-- char 0x94='\x94
--   =>	"00000000",	-- ........
 592 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........
 593 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 594 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 595 =>	"00000000",	-- ........

-- char 0x95='\x95
--   =>	"00000000",	-- ........
 596 =>	"11100000",	-- ###.....
--   =>	"00000000",	-- ........
 597 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 598 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 599 =>	"00000000",	-- ........

-- char 0x96='\x96
--   =>	"01111000",	-- .####...
 600 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........
 601 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 602 =>	"11001100",	-- ##..##..
--   =>	"01111110",	-- .######.
 603 =>	"00000000",	-- ........

-- char 0x97='\x97
--   =>	"00000000",	-- ........
 604 =>	"11100000",	-- ###.....
--   =>	"00000000",	-- ........
 605 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 606 =>	"11001100",	-- ##..##..
--   =>	"01111110",	-- .######.
 607 =>	"00000000",	-- ........

-- char 0x98='\x98
--   =>	"00000000",	-- ........
 608 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........
 609 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 610 =>	"01111100",	-- .#####..
--   =>	"00001100",	-- ....##..
 611 =>	"11111000",	-- #####...

-- char 0x99='\x99
--   =>	"11000011",	-- ##....##
 612 =>	"00011000",	-- ...##...
--   =>	"00111100",	-- ..####..
 613 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 614 =>	"00111100",	-- ..####..
--   =>	"00011000",	-- ...##...
 615 =>	"00000000",	-- ........

-- char 0x9a='\x9a
--   =>	"11001100",	-- ##..##..
 616 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 617 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 618 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 619 =>	"00000000",	-- ........

-- char 0x9b='\x9b
--   =>	"00011000",	-- ...##...
 620 =>	"00011000",	-- ...##...
--   =>	"01111110",	-- .######.
 621 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 622 =>	"01111110",	-- .######.
--   =>	"00011000",	-- ...##...
 623 =>	"00011000",	-- ...##...

-- char 0x9c='\x9c
--   =>	"00111000",	-- ..###...
 624 =>	"01101100",	-- .##.##..
--   =>	"01100100",	-- .##..#..
 625 =>	"11110000",	-- ####....
--   =>	"01100000",	-- .##.....
 626 =>	"11100110",	-- ###..##.
--   =>	"11111100",	-- ######..
 627 =>	"00000000",	-- ........

-- char 0x9d='\x9d
--   =>	"11001100",	-- ##..##..
 628 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 629 =>	"11111100",	-- ######..
--   =>	"00110000",	-- ..##....
 630 =>	"11111100",	-- ######..
--   =>	"00110000",	-- ..##....
 631 =>	"00110000",	-- ..##....

-- char 0x9e='\x9e
--   =>	"11111000",	-- #####...
 632 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 633 =>	"11111010",	-- #####.#.
--   =>	"11000110",	-- ##...##.
 634 =>	"11001111",	-- ##..####
--   =>	"11000110",	-- ##...##.
 635 =>	"11000111",	-- ##...###

-- char 0x9f='\x9f
--   =>	"00001110",	-- ....###.
 636 =>	"00011011",	-- ...##.##
--   =>	"00011000",	-- ...##...
 637 =>	"00111100",	-- ..####..
--   =>	"00011000",	-- ...##...
 638 =>	"00011000",	-- ...##...
--   =>	"11011000",	-- ##.##...
 639 =>	"01110000",	-- .###....

-- char 0xa0='\xa0
--   =>	"00011100",	-- ...###..
 640 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 641 =>	"00001100",	-- ....##..
--   =>	"01111100",	-- .#####..
 642 =>	"11001100",	-- ##..##..
--   =>	"01111110",	-- .######.
 643 =>	"00000000",	-- ........

-- char 0xa1='\xa1
--   =>	"00111000",	-- ..###...
 644 =>	"00000000",	-- ........
--   =>	"01110000",	-- .###....
 645 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 646 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 647 =>	"00000000",	-- ........

-- char 0xa2='\xa2
--   =>	"00000000",	-- ........
 648 =>	"00011100",	-- ...###..
--   =>	"00000000",	-- ........
 649 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 650 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 651 =>	"00000000",	-- ........

-- char 0xa3='\xa3
--   =>	"00000000",	-- ........
 652 =>	"00011100",	-- ...###..
--   =>	"00000000",	-- ........
 653 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 654 =>	"11001100",	-- ##..##..
--   =>	"01111110",	-- .######.
 655 =>	"00000000",	-- ........

-- char 0xa4='\xa4
--   =>	"00000000",	-- ........
 656 =>	"11111000",	-- #####...
--   =>	"00000000",	-- ........
 657 =>	"11111000",	-- #####...
--   =>	"11001100",	-- ##..##..
 658 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 659 =>	"00000000",	-- ........

-- char 0xa5='\xa5
--   =>	"11111100",	-- ######..
 660 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 661 =>	"11101100",	-- ###.##..
--   =>	"11111100",	-- ######..
 662 =>	"11011100",	-- ##.###..
--   =>	"11001100",	-- ##..##..
 663 =>	"00000000",	-- ........

-- char 0xa6='\xa6
--   =>	"00111100",	-- ..####..
 664 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 665 =>	"00111110",	-- ..#####.
--   =>	"00000000",	-- ........
 666 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........
 667 =>	"00000000",	-- ........

-- char 0xa7='\xa7
--   =>	"00111000",	-- ..###...
 668 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 669 =>	"00111000",	-- ..###...
--   =>	"00000000",	-- ........
 670 =>	"01111100",	-- .#####..
--   =>	"00000000",	-- ........
 671 =>	"00000000",	-- ........

-- char 0xa8='\xa8
--   =>	"00110000",	-- ..##....
 672 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 673 =>	"01100000",	-- .##.....
--   =>	"11000000",	-- ##......
 674 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 675 =>	"00000000",	-- ........

-- char 0xa9='\xa9
--   =>	"00000000",	-- ........
 676 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 677 =>	"11111100",	-- ######..
--   =>	"11000000",	-- ##......
 678 =>	"11000000",	-- ##......
--   =>	"00000000",	-- ........
 679 =>	"00000000",	-- ........

-- char 0xaa='\xaa
--   =>	"00000000",	-- ........
 680 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 681 =>	"11111100",	-- ######..
--   =>	"00001100",	-- ....##..
 682 =>	"00001100",	-- ....##..
--   =>	"00000000",	-- ........
 683 =>	"00000000",	-- ........

-- char 0xab='\xab
--   =>	"11000011",	-- ##....##
 684 =>	"11000110",	-- ##...##.
--   =>	"11001100",	-- ##..##..
 685 =>	"11011110",	-- ##.####.
--   =>	"00110011",	-- ..##..##
 686 =>	"01100110",	-- .##..##.
--   =>	"11001100",	-- ##..##..
 687 =>	"00001111",	-- ....####

-- char 0xac='\xac
--   =>	"11000011",	-- ##....##
 688 =>	"11000110",	-- ##...##.
--   =>	"11001100",	-- ##..##..
 689 =>	"11011011",	-- ##.##.##
--   =>	"00110111",	-- ..##.###
 690 =>	"01101111",	-- .##.####
--   =>	"11001111",	-- ##..####
 691 =>	"00000011",	-- ......##

-- char 0xad='\xad
--   =>	"00011000",	-- ...##...
 692 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........
 693 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 694 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 695 =>	"00000000",	-- ........

-- char 0xae='\xae
--   =>	"00000000",	-- ........
 696 =>	"00110011",	-- ..##..##
--   =>	"01100110",	-- .##..##.
 697 =>	"11001100",	-- ##..##..
--   =>	"01100110",	-- .##..##.
 698 =>	"00110011",	-- ..##..##
--   =>	"00000000",	-- ........
 699 =>	"00000000",	-- ........

-- char 0xaf='\xaf
--   =>	"00000000",	-- ........
 700 =>	"11001100",	-- ##..##..
--   =>	"01100110",	-- .##..##.
 701 =>	"00110011",	-- ..##..##
--   =>	"01100110",	-- .##..##.
 702 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........
 703 =>	"00000000",	-- ........

-- char 0xb0='\xb0
--   =>	"00100010",	-- ..#...#.
 704 =>	"10001000",	-- #...#...
--   =>	"00100010",	-- ..#...#.
 705 =>	"10001000",	-- #...#...
--   =>	"00100010",	-- ..#...#.
 706 =>	"10001000",	-- #...#...
--   =>	"00100010",	-- ..#...#.
 707 =>	"10001000",	-- #...#...

-- char 0xb1='\xb1
--   =>	"01010101",	-- .#.#.#.#
 708 =>	"10101010",	-- #.#.#.#.
--   =>	"01010101",	-- .#.#.#.#
 709 =>	"10101010",	-- #.#.#.#.
--   =>	"01010101",	-- .#.#.#.#
 710 =>	"10101010",	-- #.#.#.#.
--   =>	"01010101",	-- .#.#.#.#
 711 =>	"10101010",	-- #.#.#.#.

-- char 0xb2='\xb2
--   =>	"11011011",	-- ##.##.##
 712 =>	"01110111",	-- .###.###
--   =>	"11011011",	-- ##.##.##
 713 =>	"11101110",	-- ###.###.
--   =>	"11011011",	-- ##.##.##
 714 =>	"01110111",	-- .###.###
--   =>	"11011011",	-- ##.##.##
 715 =>	"11101110",	-- ###.###.

-- char 0xb3='\xb3
--   =>	"00011000",	-- ...##...
 716 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 717 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 718 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 719 =>	"00011000",	-- ...##...

-- char 0xb4='\xb4
--   =>	"00011000",	-- ...##...
 720 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 721 =>	"00011000",	-- ...##...
--   =>	"11111000",	-- #####...
 722 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 723 =>	"00011000",	-- ...##...

-- char 0xb5='\xb5
--   =>	"00011000",	-- ...##...
 724 =>	"00011000",	-- ...##...
--   =>	"11111000",	-- #####...
 725 =>	"00011000",	-- ...##...
--   =>	"11111000",	-- #####...
 726 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 727 =>	"00011000",	-- ...##...

-- char 0xb6='\xb6
--   =>	"00110110",	-- ..##.##.
 728 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 729 =>	"00110110",	-- ..##.##.
--   =>	"11110110",	-- ####.##.
 730 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 731 =>	"00110110",	-- ..##.##.

-- char 0xb7='\xb7
--   =>	"00000000",	-- ........
 732 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 733 =>	"00000000",	-- ........
--   =>	"11111110",	-- #######.
 734 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 735 =>	"00110110",	-- ..##.##.

-- char 0xb8='\xb8
--   =>	"00000000",	-- ........
 736 =>	"00000000",	-- ........
--   =>	"11111000",	-- #####...
 737 =>	"00011000",	-- ...##...
--   =>	"11111000",	-- #####...
 738 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 739 =>	"00011000",	-- ...##...

-- char 0xb9='\xb9
--   =>	"00110110",	-- ..##.##.
 740 =>	"00110110",	-- ..##.##.
--   =>	"11110110",	-- ####.##.
 741 =>	"00000110",	-- .....##.
--   =>	"11110110",	-- ####.##.
 742 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 743 =>	"00110110",	-- ..##.##.

-- char 0xba='\xba
--   =>	"00110110",	-- ..##.##.
 744 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 745 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 746 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 747 =>	"00110110",	-- ..##.##.

-- char 0xbb='\xbb
--   =>	"00000000",	-- ........
 748 =>	"00000000",	-- ........
--   =>	"11111110",	-- #######.
 749 =>	"00000110",	-- .....##.
--   =>	"11110110",	-- ####.##.
 750 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 751 =>	"00110110",	-- ..##.##.

-- char 0xbc='\xbc
--   =>	"00110110",	-- ..##.##.
 752 =>	"00110110",	-- ..##.##.
--   =>	"11110110",	-- ####.##.
 753 =>	"00000110",	-- .....##.
--   =>	"11111110",	-- #######.
 754 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 755 =>	"00000000",	-- ........

-- char 0xbd='\xbd
--   =>	"00110110",	-- ..##.##.
 756 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 757 =>	"00110110",	-- ..##.##.
--   =>	"11111110",	-- #######.
 758 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 759 =>	"00000000",	-- ........

-- char 0xbe='\xbe
--   =>	"00011000",	-- ...##...
 760 =>	"00011000",	-- ...##...
--   =>	"11111000",	-- #####...
 761 =>	"00011000",	-- ...##...
--   =>	"11111000",	-- #####...
 762 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 763 =>	"00000000",	-- ........

-- char 0xbf='\xbf
--   =>	"00000000",	-- ........
 764 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 765 =>	"00000000",	-- ........
--   =>	"11111000",	-- #####...
 766 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 767 =>	"00011000",	-- ...##...

-- char 0xc0='\xc0
--   =>	"00011000",	-- ...##...
 768 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 769 =>	"00011000",	-- ...##...
--   =>	"00011111",	-- ...#####
 770 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 771 =>	"00000000",	-- ........

-- char 0xc1='\xc1
--   =>	"00011000",	-- ...##...
 772 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 773 =>	"00011000",	-- ...##...
--   =>	"11111111",	-- ########
 774 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 775 =>	"00000000",	-- ........

-- char 0xc2='\xc2
--   =>	"00000000",	-- ........
 776 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 777 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 778 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 779 =>	"00011000",	-- ...##...

-- char 0xc3='\xc3
--   =>	"00011000",	-- ...##...
 780 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 781 =>	"00011000",	-- ...##...
--   =>	"00011111",	-- ...#####
 782 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 783 =>	"00011000",	-- ...##...

-- char 0xc4='\xc4
--   =>	"00000000",	-- ........
 784 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 785 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 786 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 787 =>	"00000000",	-- ........

-- char 0xc5='\xc5
--   =>	"00011000",	-- ...##...
 788 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 789 =>	"00011000",	-- ...##...
--   =>	"11111111",	-- ########
 790 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 791 =>	"00011000",	-- ...##...

-- char 0xc6='\xc6
--   =>	"00011000",	-- ...##...
 792 =>	"00011000",	-- ...##...
--   =>	"00011111",	-- ...#####
 793 =>	"00011000",	-- ...##...
--   =>	"00011111",	-- ...#####
 794 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 795 =>	"00011000",	-- ...##...

-- char 0xc7='\xc7
--   =>	"00110110",	-- ..##.##.
 796 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 797 =>	"00110110",	-- ..##.##.
--   =>	"00110111",	-- ..##.###
 798 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 799 =>	"00110110",	-- ..##.##.

-- char 0xc8='\xc8
--   =>	"00110110",	-- ..##.##.
 800 =>	"00110110",	-- ..##.##.
--   =>	"00110111",	-- ..##.###
 801 =>	"00110000",	-- ..##....
--   =>	"00111111",	-- ..######
 802 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 803 =>	"00000000",	-- ........

-- char 0xc9='\xc9
--   =>	"00000000",	-- ........
 804 =>	"00000000",	-- ........
--   =>	"00111111",	-- ..######
 805 =>	"00110000",	-- ..##....
--   =>	"00110111",	-- ..##.###
 806 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 807 =>	"00110110",	-- ..##.##.

-- char 0xca='\xca
--   =>	"00110110",	-- ..##.##.
 808 =>	"00110110",	-- ..##.##.
--   =>	"11110111",	-- ####.###
 809 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 810 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 811 =>	"00000000",	-- ........

-- char 0xcb='\xcb
--   =>	"00000000",	-- ........
 812 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 813 =>	"00000000",	-- ........
--   =>	"11110111",	-- ####.###
 814 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 815 =>	"00110110",	-- ..##.##.

-- char 0xcc='\xcc
--   =>	"00110110",	-- ..##.##.
 816 =>	"00110110",	-- ..##.##.
--   =>	"00110111",	-- ..##.###
 817 =>	"00110000",	-- ..##....
--   =>	"00110111",	-- ..##.###
 818 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 819 =>	"00110110",	-- ..##.##.

-- char 0xcd='\xcd
--   =>	"00000000",	-- ........
 820 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 821 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 822 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 823 =>	"00000000",	-- ........

-- char 0xce='\xce
--   =>	"00110110",	-- ..##.##.
 824 =>	"00110110",	-- ..##.##.
--   =>	"11110111",	-- ####.###
 825 =>	"00000000",	-- ........
--   =>	"11110111",	-- ####.###
 826 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 827 =>	"00110110",	-- ..##.##.

-- char 0xcf='\xcf
--   =>	"00011000",	-- ...##...
 828 =>	"00011000",	-- ...##...
--   =>	"11111111",	-- ########
 829 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 830 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 831 =>	"00000000",	-- ........

-- char 0xd0='\xd0
--   =>	"00110110",	-- ..##.##.
 832 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 833 =>	"00110110",	-- ..##.##.
--   =>	"11111111",	-- ########
 834 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 835 =>	"00000000",	-- ........

-- char 0xd1='\xd1
--   =>	"00000000",	-- ........
 836 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 837 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 838 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 839 =>	"00011000",	-- ...##...

-- char 0xd2='\xd2
--   =>	"00000000",	-- ........
 840 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 841 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 842 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 843 =>	"00110110",	-- ..##.##.

-- char 0xd3='\xd3
--   =>	"00110110",	-- ..##.##.
 844 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 845 =>	"00110110",	-- ..##.##.
--   =>	"00111111",	-- ..######
 846 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 847 =>	"00000000",	-- ........

-- char 0xd4='\xd4
--   =>	"00011000",	-- ...##...
 848 =>	"00011000",	-- ...##...
--   =>	"00011111",	-- ...#####
 849 =>	"00011000",	-- ...##...
--   =>	"00011111",	-- ...#####
 850 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 851 =>	"00000000",	-- ........

-- char 0xd5='\xd5
--   =>	"00000000",	-- ........
 852 =>	"00000000",	-- ........
--   =>	"00011111",	-- ...#####
 853 =>	"00011000",	-- ...##...
--   =>	"00011111",	-- ...#####
 854 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 855 =>	"00011000",	-- ...##...

-- char 0xd6='\xd6
--   =>	"00000000",	-- ........
 856 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 857 =>	"00000000",	-- ........
--   =>	"00111111",	-- ..######
 858 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 859 =>	"00110110",	-- ..##.##.

-- char 0xd7='\xd7
--   =>	"00110110",	-- ..##.##.
 860 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 861 =>	"00110110",	-- ..##.##.
--   =>	"11111111",	-- ########
 862 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 863 =>	"00110110",	-- ..##.##.

-- char 0xd8='\xd8
--   =>	"00011000",	-- ...##...
 864 =>	"00011000",	-- ...##...
--   =>	"11111111",	-- ########
 865 =>	"00011000",	-- ...##...
--   =>	"11111111",	-- ########
 866 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 867 =>	"00011000",	-- ...##...

-- char 0xd9='\xd9
--   =>	"00011000",	-- ...##...
 868 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 869 =>	"00011000",	-- ...##...
--   =>	"11111000",	-- #####...
 870 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 871 =>	"00000000",	-- ........

-- char 0xda='\xda
--   =>	"00000000",	-- ........
 872 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 873 =>	"00000000",	-- ........
--   =>	"00011111",	-- ...#####
 874 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 875 =>	"00011000",	-- ...##...

-- char 0xdb='\xdb
--   =>	"11111111",	-- ########
 876 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 877 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 878 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 879 =>	"11111111",	-- ########

-- char 0xdc='\xdc
--   =>	"00000000",	-- ........
 880 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 881 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 882 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 883 =>	"11111111",	-- ########

-- char 0xdd='\xdd
--   =>	"11110000",	-- ####....
 884 =>	"11110000",	-- ####....
--   =>	"11110000",	-- ####....
 885 =>	"11110000",	-- ####....
--   =>	"11110000",	-- ####....
 886 =>	"11110000",	-- ####....
--   =>	"11110000",	-- ####....
 887 =>	"11110000",	-- ####....

-- char 0xde='\xde
--   =>	"00001111",	-- ....####
 888 =>	"00001111",	-- ....####
--   =>	"00001111",	-- ....####
 889 =>	"00001111",	-- ....####
--   =>	"00001111",	-- ....####
 890 =>	"00001111",	-- ....####
--   =>	"00001111",	-- ....####
 891 =>	"00001111",	-- ....####

-- char 0xdf='\xdf
--   =>	"11111111",	-- ########
 892 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 893 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 894 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 895 =>	"00000000",	-- ........

-- char 0xe0='\xe0
--   =>	"00000000",	-- ........
 896 =>	"00000000",	-- ........
--   =>	"01110110",	-- .###.##.
 897 =>	"11011100",	-- ##.###..
--   =>	"11001000",	-- ##..#...
 898 =>	"11011100",	-- ##.###..
--   =>	"01110110",	-- .###.##.
 899 =>	"00000000",	-- ........

-- char 0xe1='\xe1
--   =>	"00000000",	-- ........
 900 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 901 =>	"11111000",	-- #####...
--   =>	"11001100",	-- ##..##..
 902 =>	"11111000",	-- #####...
--   =>	"11000000",	-- ##......
 903 =>	"11000000",	-- ##......

-- char 0xe2='\xe2
--   =>	"00000000",	-- ........
 904 =>	"11111100",	-- ######..
--   =>	"11001100",	-- ##..##..
 905 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 906 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 907 =>	"00000000",	-- ........

-- char 0xe3='\xe3
--   =>	"00000000",	-- ........
 908 =>	"11111110",	-- #######.
--   =>	"01101100",	-- .##.##..
 909 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 910 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 911 =>	"00000000",	-- ........

-- char 0xe4='\xe4
--   =>	"11111100",	-- ######..
 912 =>	"11001100",	-- ##..##..
--   =>	"01100000",	-- .##.....
 913 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
 914 =>	"11001100",	-- ##..##..
--   =>	"11111100",	-- ######..
 915 =>	"00000000",	-- ........

-- char 0xe5='\xe5
--   =>	"00000000",	-- ........
 916 =>	"00000000",	-- ........
--   =>	"01111110",	-- .######.
 917 =>	"11011000",	-- ##.##...
--   =>	"11011000",	-- ##.##...
 918 =>	"11011000",	-- ##.##...
--   =>	"01110000",	-- .###....
 919 =>	"00000000",	-- ........

-- char 0xe6='\xe6
--   =>	"00000000",	-- ........
 920 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 921 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 922 =>	"01111100",	-- .#####..
--   =>	"01100000",	-- .##.....
 923 =>	"11000000",	-- ##......

-- char 0xe7='\xe7
--   =>	"00000000",	-- ........
 924 =>	"01110110",	-- .###.##.
--   =>	"11011100",	-- ##.###..
 925 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 926 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 927 =>	"00000000",	-- ........

-- char 0xe8='\xe8
--   =>	"11111100",	-- ######..
 928 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 929 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 930 =>	"01111000",	-- .####...
--   =>	"00110000",	-- ..##....
 931 =>	"11111100",	-- ######..

-- char 0xe9='\xe9
--   =>	"00111000",	-- ..###...
 932 =>	"01101100",	-- .##.##..
--   =>	"11000110",	-- ##...##.
 933 =>	"11111110",	-- #######.
--   =>	"11000110",	-- ##...##.
 934 =>	"01101100",	-- .##.##..
--   =>	"00111000",	-- ..###...
 935 =>	"00000000",	-- ........

-- char 0xea='\xea
--   =>	"00111000",	-- ..###...
 936 =>	"01101100",	-- .##.##..
--   =>	"11000110",	-- ##...##.
 937 =>	"11000110",	-- ##...##.
--   =>	"01101100",	-- .##.##..
 938 =>	"01101100",	-- .##.##..
--   =>	"11101110",	-- ###.###.
 939 =>	"00000000",	-- ........

-- char 0xeb='\xeb
--   =>	"00011100",	-- ...###..
 940 =>	"00110000",	-- ..##....
--   =>	"00011000",	-- ...##...
 941 =>	"01111100",	-- .#####..
--   =>	"11001100",	-- ##..##..
 942 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 943 =>	"00000000",	-- ........

-- char 0xec='\xec
--   =>	"00000000",	-- ........
 944 =>	"00000000",	-- ........
--   =>	"01111110",	-- .######.
 945 =>	"11011011",	-- ##.##.##
--   =>	"11011011",	-- ##.##.##
 946 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........
 947 =>	"00000000",	-- ........

-- char 0xed='\xed
--   =>	"00000110",	-- .....##.
 948 =>	"00001100",	-- ....##..
--   =>	"01111110",	-- .######.
 949 =>	"11011011",	-- ##.##.##
--   =>	"11011011",	-- ##.##.##
 950 =>	"01111110",	-- .######.
--   =>	"01100000",	-- .##.....
 951 =>	"11000000",	-- ##......

-- char 0xee='\xee
--   =>	"00111000",	-- ..###...
 952 =>	"01100000",	-- .##.....
--   =>	"11000000",	-- ##......
 953 =>	"11111000",	-- #####...
--   =>	"11000000",	-- ##......
 954 =>	"01100000",	-- .##.....
--   =>	"00111000",	-- ..###...
 955 =>	"00000000",	-- ........

-- char 0xef='\xef
--   =>	"01111000",	-- .####...
 956 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 957 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 958 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 959 =>	"00000000",	-- ........

-- char 0xf0='\xf0
--   =>	"00000000",	-- ........
 960 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........
 961 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........
 962 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........
 963 =>	"00000000",	-- ........

-- char 0xf1='\xf1
--   =>	"00110000",	-- ..##....
 964 =>	"00110000",	-- ..##....
--   =>	"11111100",	-- ######..
 965 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 966 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 967 =>	"00000000",	-- ........

-- char 0xf2='\xf2
--   =>	"01100000",	-- .##.....
 968 =>	"00110000",	-- ..##....
--   =>	"00011000",	-- ...##...
 969 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
 970 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 971 =>	"00000000",	-- ........

-- char 0xf3='\xf3
--   =>	"00011000",	-- ...##...
 972 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
 973 =>	"00110000",	-- ..##....
--   =>	"00011000",	-- ...##...
 974 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 975 =>	"00000000",	-- ........

-- char 0xf4='\xf4
--   =>	"00001110",	-- ....###.
 976 =>	"00011011",	-- ...##.##
--   =>	"00011011",	-- ...##.##
 977 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 978 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 979 =>	"00011000",	-- ...##...

-- char 0xf5='\xf5
--   =>	"00011000",	-- ...##...
 980 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 981 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 982 =>	"11011000",	-- ##.##...
--   =>	"11011000",	-- ##.##...
 983 =>	"01110000",	-- .###....

-- char 0xf6='\xf6
--   =>	"00110000",	-- ..##....
 984 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 985 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........
 986 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 987 =>	"00000000",	-- ........

-- char 0xf7='\xf7
--   =>	"00000000",	-- ........
 988 =>	"01110110",	-- .###.##.
--   =>	"11011100",	-- ##.###..
 989 =>	"00000000",	-- ........
--   =>	"01110110",	-- .###.##.
 990 =>	"11011100",	-- ##.###..
--   =>	"00000000",	-- ........
 991 =>	"00000000",	-- ........

-- char 0xf8='\xf8
--   =>	"00111000",	-- ..###...
 992 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 993 =>	"00111000",	-- ..###...
--   =>	"00000000",	-- ........
 994 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 995 =>	"00000000",	-- ........

-- char 0xf9='\xf9
--   =>	"00000000",	-- ........
 996 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 997 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 998 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 999 =>	"00000000",	-- ........

-- char 0xfa='\xfa
--   =>	"00000000",	-- ........
1000 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1001 =>	"00000000",	-- ........
--   =>	"00011000",	-- ...##...
1002 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1003 =>	"00000000",	-- ........

-- char 0xfb='\xfb
--   =>	"00001111",	-- ....####
1004 =>	"00001100",	-- ....##..
--   =>	"00001100",	-- ....##..
1005 =>	"00001100",	-- ....##..
--   =>	"11101100",	-- ###.##..
1006 =>	"01101100",	-- .##.##..
--   =>	"00111100",	-- ..####..
1007 =>	"00011100",	-- ...###..

-- char 0xfc='\xfc
--   =>	"01111000",	-- .####...
1008 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
1009 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
1010 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1011 =>	"00000000",	-- ........

-- char 0xfd='\xfd
--   =>	"01110000",	-- .###....
1012 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
1013 =>	"01100000",	-- .##.....
--   =>	"01111000",	-- .####...
1014 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1015 =>	"00000000",	-- ........

-- char 0xfe='\xfe
--   =>	"00000000",	-- ........
1016 =>	"00000000",	-- ........
--   =>	"00111100",	-- ..####..
1017 =>	"00111100",	-- ..####..
--   =>	"00111100",	-- ..####..
1018 =>	"00111100",	-- ..####..
--   =>	"00000000",	-- ........
1019 =>	"00000000",	-- ........

-- char 0xff='\xff
--   =>	"00000000",	-- ........
1020 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1021 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1022 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1023 =>	"00000000"	-- ........
);
	attribute syn_ramstyle: string;
	attribute syn_ramstyle of mem: signal is "no_rw_check";
begin
	process (clka_i) -- Using port a.
	begin
	if (rising_edge(clka_i)) then
		if (wea_i = '1') then
		mem(conv_integer(addra_i)) <= dina_i;
			-- Using address bus a.
		end if;
		douta_o <= mem(conv_integer(addra_i));
	end if;
	end process;
	process (clkb_i) -- Using port b.
	begin
	if (rising_edge(clkb_i)) then
		if (web_i = '1') then
		mem(conv_integer(addrb_i)) <= dinb_i;
			-- Using address bus b.
		end if;
		doutb_o <= mem(conv_integer(addrb_i));
	end if;
	end process;
end rtl;
