library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
  
entity Sweet32_SRAM_upper is

   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      addr_i  : in  std_logic_vector(11 downto 0);
      write_i : in  std_logic_vector(7 downto 0);
      read_o  : out std_logic_vector(7 downto 0)
	);
end entity Sweet32_SRAM_upper;

architecture behavioral of Sweet32_SRAM_upper is
   type ram_type is array(4095 downto 0) of std_logic_vector(7 downto 0);
   signal addr_r  : std_logic_vector(11 downto 0);

   signal ram : ram_type :=
(
 
 -- Test program, upper byte (MSB) of 16-bit (byte-addressable) ROM

   0 => x"90",
   1 => x"60",
   2 => x"00",
   3 => x"00",
   4 => x"B0",
   5 => x"0E",
   6 => x"1E",
   7 => x"E0",
   8 => x"AE",
   9 => x"E1",
  10 => x"AE",
  11 => x"E2",
  12 => x"AE",
  13 => x"E3",
  14 => x"AE",
  15 => x"E4",
  16 => x"AE",
  17 => x"E5",
  18 => x"AE",
  19 => x"E6",
  20 => x"AE",
  21 => x"E7",
  22 => x"AE",
  23 => x"E8",
  24 => x"AE",
  25 => x"E9",
  26 => x"AE",
  27 => x"EA",
  28 => x"AE",
  29 => x"EB",
  30 => x"AE",
  31 => x"EC",
  32 => x"AE",
  33 => x"ED",
  34 => x"AE",
  35 => x"B0",
  36 => x"0F",
  37 => x"10",
  38 => x"E0",
  39 => x"AE",
  40 => x"EF",
  41 => x"A0",
  42 => x"B1",
  43 => x"00",
  44 => x"70",
  45 => x"73",
  46 => x"1C",
  47 => x"70",
  48 => x"E0",
  49 => x"60",
  50 => x"B0",
  51 => x"0C",
  52 => x"B0",
  53 => x"0E",
  54 => x"16",
  55 => x"F1",
  56 => x"B0",
  57 => x"0C",
  58 => x"90",
  59 => x"64",
  60 => x"73",
  61 => x"1C",
  62 => x"70",
  63 => x"E0",
  64 => x"B0",
  65 => x"0F",
  66 => x"1E",
  67 => x"B0",
  68 => x"0E",
  69 => x"1F",
  70 => x"F1",
  71 => x"F1",
  72 => x"AF",
  73 => x"F1",
  74 => x"AF",
  75 => x"F1",
  76 => x"AF",
  77 => x"F1",
  78 => x"AF",
  79 => x"F1",
  80 => x"AF",
  81 => x"F1",
  82 => x"AF",
  83 => x"F1",
  84 => x"AF",
  85 => x"F1",
  86 => x"AF",
  87 => x"F1",
  88 => x"AF",
  89 => x"F1",
  90 => x"AF",
  91 => x"F1",
  92 => x"AF",
  93 => x"F1",
  94 => x"AF",
  95 => x"F1",
  96 => x"9A",
  97 => x"C3",
  98 => x"B0",
  99 => x"0F",
 100 => x"11",
 101 => x"7F",
 102 => x"11",
 103 => x"C2",
 104 => x"01",
 105 => x"B0",
 106 => x"0E",
 107 => x"10",
 108 => x"E1",
 109 => x"B0",
 110 => x"0E",
 111 => x"10",
 112 => x"E1",
 113 => x"B0",
 114 => x"0A",
 115 => x"90",
 116 => x"64",
 117 => x"AD",
 118 => x"B0",
 119 => x"0E",
 120 => x"16",
 121 => x"F0",
 122 => x"D0",
 123 => x"A6",
 124 => x"B0",
 125 => x"FF",
 126 => x"F0",
 127 => x"A5",
 128 => x"90",
 129 => x"63",
 130 => x"A2",
 131 => x"A6",
 132 => x"36",
 133 => x"6F",
 134 => x"23",
 135 => x"30",
 136 => x"60",
 137 => x"90",
 138 => x"64",
 139 => x"72",
 140 => x"90",
 141 => x"64",
 142 => x"A7",
 143 => x"90",
 144 => x"64",
 145 => x"B0",
 146 => x"0C",
 147 => x"90",
 148 => x"64",
 149 => x"B0",
 150 => x"0B",
 151 => x"90",
 152 => x"64",
 153 => x"90",
 154 => x"64",
 155 => x"9F",
 156 => x"74",
 157 => x"22",
 158 => x"30",
 159 => x"62",
 160 => x"74",
 161 => x"22",
 162 => x"30",
 163 => x"60",
 164 => x"74",
 165 => x"22",
 166 => x"30",
 167 => x"60",
 168 => x"74",
 169 => x"22",
 170 => x"30",
 171 => x"62",
 172 => x"75",
 173 => x"22",
 174 => x"30",
 175 => x"62",
 176 => x"75",
 177 => x"22",
 178 => x"30",
 179 => x"63",
 180 => x"74",
 181 => x"22",
 182 => x"30",
 183 => x"60",
 184 => x"75",
 185 => x"22",
 186 => x"30",
 187 => x"63",
 188 => x"70",
 189 => x"22",
 190 => x"30",
 191 => x"60",
 192 => x"B0",
 193 => x"0B",
 194 => x"64",
 195 => x"AE",
 196 => x"EF",
 197 => x"B0",
 198 => x"0B",
 199 => x"90",
 200 => x"64",
 201 => x"B0",
 202 => x"0E",
 203 => x"19",
 204 => x"F1",
 205 => x"70",
 206 => x"90",
 207 => x"63",
 208 => x"34",
 209 => x"60",
 210 => x"A2",
 211 => x"60",
 212 => x"AE",
 213 => x"EF",
 214 => x"B0",
 215 => x"0E",
 216 => x"19",
 217 => x"F1",
 218 => x"78",
 219 => x"16",
 220 => x"70",
 221 => x"B0",
 222 => x"0C",
 223 => x"A6",
 224 => x"B0",
 225 => x"0C",
 226 => x"90",
 227 => x"64",
 228 => x"F3",
 229 => x"A6",
 230 => x"A8",
 231 => x"90",
 232 => x"64",
 233 => x"26",
 234 => x"30",
 235 => x"60",
 236 => x"72",
 237 => x"90",
 238 => x"64",
 239 => x"70",
 240 => x"38",
 241 => x"6F",
 242 => x"6F",
 243 => x"B0",
 244 => x"0E",
 245 => x"19",
 246 => x"E6",
 247 => x"F1",
 248 => x"AE",
 249 => x"C3",
 250 => x"AE",
 251 => x"EF",
 252 => x"B0",
 253 => x"0B",
 254 => x"90",
 255 => x"64",
 256 => x"B0",
 257 => x"0E",
 258 => x"19",
 259 => x"F1",
 260 => x"70",
 261 => x"90",
 262 => x"63",
 263 => x"34",
 264 => x"60",
 265 => x"A2",
 266 => x"B0",
 267 => x"0C",
 268 => x"A6",
 269 => x"B0",
 270 => x"0C",
 271 => x"90",
 272 => x"64",
 273 => x"F3",
 274 => x"90",
 275 => x"63",
 276 => x"73",
 277 => x"90",
 278 => x"64",
 279 => x"F3",
 280 => x"70",
 281 => x"90",
 282 => x"63",
 283 => x"34",
 284 => x"60",
 285 => x"E2",
 286 => x"A6",
 287 => x"E6",
 288 => x"6F",
 289 => x"F1",
 290 => x"AE",
 291 => x"C3",
 292 => x"AE",
 293 => x"EF",
 294 => x"B0",
 295 => x"0B",
 296 => x"90",
 297 => x"64",
 298 => x"B0",
 299 => x"0E",
 300 => x"19",
 301 => x"F1",
 302 => x"70",
 303 => x"90",
 304 => x"63",
 305 => x"33",
 306 => x"61",
 307 => x"A2",
 308 => x"60",
 309 => x"AE",
 310 => x"EF",
 311 => x"B0",
 312 => x"0E",
 313 => x"19",
 314 => x"F1",
 315 => x"72",
 316 => x"16",
 317 => x"B0",
 318 => x"0C",
 319 => x"A6",
 320 => x"B0",
 321 => x"0C",
 322 => x"90",
 323 => x"63",
 324 => x"B0",
 325 => x"0C",
 326 => x"18",
 327 => x"F0",
 328 => x"F0",
 329 => x"03",
 330 => x"A8",
 331 => x"F0",
 332 => x"20",
 333 => x"30",
 334 => x"60",
 335 => x"A8",
 336 => x"A8",
 337 => x"6F",
 338 => x"F0",
 339 => x"90",
 340 => x"63",
 341 => x"72",
 342 => x"90",
 343 => x"63",
 344 => x"A8",
 345 => x"F3",
 346 => x"34",
 347 => x"60",
 348 => x"B0",
 349 => x"0C",
 350 => x"91",
 351 => x"63",
 352 => x"A6",
 353 => x"F0",
 354 => x"90",
 355 => x"63",
 356 => x"F3",
 357 => x"34",
 358 => x"60",
 359 => x"B0",
 360 => x"0C",
 361 => x"90",
 362 => x"63",
 363 => x"A6",
 364 => x"F0",
 365 => x"90",
 366 => x"63",
 367 => x"72",
 368 => x"90",
 369 => x"63",
 370 => x"A8",
 371 => x"A8",
 372 => x"70",
 373 => x"90",
 374 => x"63",
 375 => x"B0",
 376 => x"0C",
 377 => x"90",
 378 => x"63",
 379 => x"A8",
 380 => x"F3",
 381 => x"F0",
 382 => x"A6",
 383 => x"70",
 384 => x"41",
 385 => x"60",
 386 => x"61",
 387 => x"41",
 388 => x"60",
 389 => x"70",
 390 => x"03",
 391 => x"90",
 392 => x"62",
 393 => x"61",
 394 => x"41",
 395 => x"60",
 396 => x"7F",
 397 => x"03",
 398 => x"D0",
 399 => x"D0",
 400 => x"D0",
 401 => x"D0",
 402 => x"90",
 403 => x"62",
 404 => x"61",
 405 => x"41",
 406 => x"60",
 407 => x"B0",
 408 => x"0F",
 409 => x"03",
 410 => x"33",
 411 => x"60",
 412 => x"C2",
 413 => x"13",
 414 => x"13",
 415 => x"13",
 416 => x"90",
 417 => x"63",
 418 => x"61",
 419 => x"41",
 420 => x"60",
 421 => x"B0",
 422 => x"0F",
 423 => x"03",
 424 => x"C1",
 425 => x"A4",
 426 => x"F0",
 427 => x"13",
 428 => x"33",
 429 => x"60",
 430 => x"B1",
 431 => x"00",
 432 => x"F0",
 433 => x"13",
 434 => x"13",
 435 => x"13",
 436 => x"A3",
 437 => x"90",
 438 => x"63",
 439 => x"60",
 440 => x"41",
 441 => x"60",
 442 => x"F0",
 443 => x"70",
 444 => x"03",
 445 => x"90",
 446 => x"62",
 447 => x"72",
 448 => x"90",
 449 => x"63",
 450 => x"F0",
 451 => x"70",
 452 => x"C0",
 453 => x"03",
 454 => x"90",
 455 => x"62",
 456 => x"60",
 457 => x"41",
 458 => x"60",
 459 => x"70",
 460 => x"C0",
 461 => x"03",
 462 => x"90",
 463 => x"62",
 464 => x"B0",
 465 => x"0C",
 466 => x"90",
 467 => x"63",
 468 => x"F0",
 469 => x"71",
 470 => x"03",
 471 => x"90",
 472 => x"63",
 473 => x"60",
 474 => x"41",
 475 => x"60",
 476 => x"7F",
 477 => x"03",
 478 => x"D0",
 479 => x"D0",
 480 => x"D0",
 481 => x"D0",
 482 => x"9D",
 483 => x"62",
 484 => x"41",
 485 => x"60",
 486 => x"7F",
 487 => x"03",
 488 => x"D0",
 489 => x"D0",
 490 => x"D0",
 491 => x"D0",
 492 => x"90",
 493 => x"62",
 494 => x"72",
 495 => x"90",
 496 => x"63",
 497 => x"F0",
 498 => x"70",
 499 => x"03",
 500 => x"90",
 501 => x"62",
 502 => x"60",
 503 => x"41",
 504 => x"60",
 505 => x"7F",
 506 => x"03",
 507 => x"D0",
 508 => x"D0",
 509 => x"D0",
 510 => x"D0",
 511 => x"90",
 512 => x"62",
 513 => x"72",
 514 => x"90",
 515 => x"63",
 516 => x"74",
 517 => x"9E",
 518 => x"63",
 519 => x"41",
 520 => x"60",
 521 => x"74",
 522 => x"9B",
 523 => x"63",
 524 => x"41",
 525 => x"60",
 526 => x"7F",
 527 => x"03",
 528 => x"D0",
 529 => x"D0",
 530 => x"D0",
 531 => x"D0",
 532 => x"90",
 533 => x"62",
 534 => x"B0",
 535 => x"0C",
 536 => x"90",
 537 => x"63",
 538 => x"F0",
 539 => x"70",
 540 => x"01",
 541 => x"B0",
 542 => x"0F",
 543 => x"01",
 544 => x"D0",
 545 => x"D0",
 546 => x"D0",
 547 => x"D0",
 548 => x"13",
 549 => x"90",
 550 => x"62",
 551 => x"60",
 552 => x"41",
 553 => x"60",
 554 => x"7F",
 555 => x"03",
 556 => x"D0",
 557 => x"D0",
 558 => x"D0",
 559 => x"D0",
 560 => x"90",
 561 => x"62",
 562 => x"72",
 563 => x"90",
 564 => x"63",
 565 => x"F0",
 566 => x"70",
 567 => x"01",
 568 => x"B0",
 569 => x"0F",
 570 => x"01",
 571 => x"D0",
 572 => x"D0",
 573 => x"D0",
 574 => x"D0",
 575 => x"13",
 576 => x"33",
 577 => x"60",
 578 => x"7F",
 579 => x"C2",
 580 => x"13",
 581 => x"13",
 582 => x"13",
 583 => x"96",
 584 => x"62",
 585 => x"41",
 586 => x"60",
 587 => x"7F",
 588 => x"03",
 589 => x"D0",
 590 => x"D0",
 591 => x"D0",
 592 => x"D0",
 593 => x"90",
 594 => x"61",
 595 => x"B0",
 596 => x"0C",
 597 => x"90",
 598 => x"62",
 599 => x"A6",
 600 => x"F0",
 601 => x"95",
 602 => x"62",
 603 => x"41",
 604 => x"60",
 605 => x"7F",
 606 => x"03",
 607 => x"D0",
 608 => x"D0",
 609 => x"D0",
 610 => x"D0",
 611 => x"90",
 612 => x"61",
 613 => x"B0",
 614 => x"0C",
 615 => x"90",
 616 => x"62",
 617 => x"A6",
 618 => x"F1",
 619 => x"94",
 620 => x"62",
 621 => x"41",
 622 => x"60",
 623 => x"7F",
 624 => x"03",
 625 => x"D0",
 626 => x"D0",
 627 => x"D0",
 628 => x"D0",
 629 => x"90",
 630 => x"61",
 631 => x"72",
 632 => x"90",
 633 => x"62",
 634 => x"F0",
 635 => x"70",
 636 => x"C0",
 637 => x"03",
 638 => x"90",
 639 => x"61",
 640 => x"6F",
 641 => x"41",
 642 => x"60",
 643 => x"7F",
 644 => x"03",
 645 => x"D0",
 646 => x"D0",
 647 => x"D0",
 648 => x"D0",
 649 => x"90",
 650 => x"61",
 651 => x"72",
 652 => x"90",
 653 => x"62",
 654 => x"6F",
 655 => x"7F",
 656 => x"03",
 657 => x"D0",
 658 => x"D0",
 659 => x"D0",
 660 => x"D0",
 661 => x"90",
 662 => x"61",
 663 => x"72",
 664 => x"90",
 665 => x"62",
 666 => x"F0",
 667 => x"70",
 668 => x"C0",
 669 => x"03",
 670 => x"90",
 671 => x"61",
 672 => x"B0",
 673 => x"0C",
 674 => x"90",
 675 => x"62",
 676 => x"F0",
 677 => x"70",
 678 => x"03",
 679 => x"33",
 680 => x"60",
 681 => x"A3",
 682 => x"72",
 683 => x"90",
 684 => x"62",
 685 => x"70",
 686 => x"C2",
 687 => x"03",
 688 => x"A3",
 689 => x"90",
 690 => x"62",
 691 => x"A8",
 692 => x"F3",
 693 => x"10",
 694 => x"16",
 695 => x"46",
 696 => x"6E",
 697 => x"B0",
 698 => x"0E",
 699 => x"19",
 700 => x"E6",
 701 => x"F1",
 702 => x"AE",
 703 => x"C3",
 704 => x"AE",
 705 => x"EF",
 706 => x"AC",
 707 => x"F0",
 708 => x"B0",
 709 => x"0B",
 710 => x"90",
 711 => x"62",
 712 => x"70",
 713 => x"B0",
 714 => x"0C",
 715 => x"90",
 716 => x"62",
 717 => x"A6",
 718 => x"90",
 719 => x"62",
 720 => x"90",
 721 => x"62",
 722 => x"90",
 723 => x"62",
 724 => x"A2",
 725 => x"AC",
 726 => x"F0",
 727 => x"36",
 728 => x"6F",
 729 => x"AC",
 730 => x"E6",
 731 => x"70",
 732 => x"90",
 733 => x"62",
 734 => x"70",
 735 => x"90",
 736 => x"62",
 737 => x"75",
 738 => x"25",
 739 => x"30",
 740 => x"6F",
 741 => x"A8",
 742 => x"38",
 743 => x"6F",
 744 => x"B0",
 745 => x"0C",
 746 => x"90",
 747 => x"62",
 748 => x"A6",
 749 => x"90",
 750 => x"62",
 751 => x"90",
 752 => x"62",
 753 => x"F1",
 754 => x"AE",
 755 => x"C3",
 756 => x"AE",
 757 => x"EF",
 758 => x"B0",
 759 => x"0B",
 760 => x"90",
 761 => x"62",
 762 => x"B0",
 763 => x"0E",
 764 => x"15",
 765 => x"F1",
 766 => x"70",
 767 => x"90",
 768 => x"61",
 769 => x"34",
 770 => x"60",
 771 => x"E2",
 772 => x"6D",
 773 => x"F1",
 774 => x"AE",
 775 => x"C3",
 776 => x"AE",
 777 => x"EF",
 778 => x"70",
 779 => x"C1",
 780 => x"70",
 781 => x"F0",
 782 => x"30",
 783 => x"60",
 784 => x"44",
 785 => x"6F",
 786 => x"B0",
 787 => x"0B",
 788 => x"90",
 789 => x"62",
 790 => x"70",
 791 => x"70",
 792 => x"90",
 793 => x"62",
 794 => x"75",
 795 => x"20",
 796 => x"30",
 797 => x"60",
 798 => x"AB",
 799 => x"6F",
 800 => x"75",
 801 => x"20",
 802 => x"30",
 803 => x"60",
 804 => x"71",
 805 => x"20",
 806 => x"30",
 807 => x"60",
 808 => x"A5",
 809 => x"70",
 810 => x"35",
 811 => x"6F",
 812 => x"60",
 813 => x"90",
 814 => x"62",
 815 => x"77",
 816 => x"20",
 817 => x"30",
 818 => x"60",
 819 => x"90",
 820 => x"60",
 821 => x"B0",
 822 => x"32",
 823 => x"20",
 824 => x"30",
 825 => x"60",
 826 => x"90",
 827 => x"60",
 828 => x"B0",
 829 => x"32",
 830 => x"20",
 831 => x"30",
 832 => x"60",
 833 => x"B0",
 834 => x"0E",
 835 => x"18",
 836 => x"90",
 837 => x"60",
 838 => x"70",
 839 => x"F0",
 840 => x"30",
 841 => x"6F",
 842 => x"E3",
 843 => x"36",
 844 => x"E6",
 845 => x"36",
 846 => x"F1",
 847 => x"90",
 848 => x"60",
 849 => x"B1",
 850 => x"FF",
 851 => x"00",
 852 => x"40",
 853 => x"60",
 854 => x"70",
 855 => x"F0",
 856 => x"30",
 857 => x"6F",
 858 => x"E3",
 859 => x"A6",
 860 => x"F1",
 861 => x"90",
 862 => x"60",
 863 => x"A2",
 864 => x"E4",
 865 => x"A8",
 866 => x"A7",
 867 => x"37",
 868 => x"60",
 869 => x"72",
 870 => x"9F",
 871 => x"61",
 872 => x"70",
 873 => x"B0",
 874 => x"0C",
 875 => x"93",
 876 => x"61",
 877 => x"90",
 878 => x"60",
 879 => x"B0",
 880 => x"64",
 881 => x"20",
 882 => x"30",
 883 => x"6F",
 884 => x"90",
 885 => x"60",
 886 => x"A2",
 887 => x"B0",
 888 => x"0B",
 889 => x"B0",
 890 => x"0E",
 891 => x"14",
 892 => x"F1",
 893 => x"70",
 894 => x"90",
 895 => x"61",
 896 => x"72",
 897 => x"90",
 898 => x"61",
 899 => x"B0",
 900 => x"0E",
 901 => x"14",
 902 => x"F1",
 903 => x"16",
 904 => x"90",
 905 => x"61",
 906 => x"B0",
 907 => x"0B",
 908 => x"90",
 909 => x"61",
 910 => x"B0",
 911 => x"0E",
 912 => x"10",
 913 => x"F1",
 914 => x"B0",
 915 => x"FF",
 916 => x"F0",
 917 => x"A5",
 918 => x"90",
 919 => x"60",
 920 => x"A2",
 921 => x"A6",
 922 => x"36",
 923 => x"6F",
 924 => x"A2",
 925 => x"A2",
 926 => x"90",
 927 => x"61",
 928 => x"B0",
 929 => x"0C",
 930 => x"90",
 931 => x"28",
 932 => x"30",
 933 => x"60",
 934 => x"B0",
 935 => x"0C",
 936 => x"9C",
 937 => x"61",
 938 => x"AB",
 939 => x"3B",
 940 => x"6C",
 941 => x"90",
 942 => x"61",
 943 => x"F1",
 944 => x"AE",
 945 => x"C3",
 946 => x"AE",
 947 => x"EF",
 948 => x"90",
 949 => x"61",
 950 => x"A2",
 951 => x"90",
 952 => x"61",
 953 => x"C0",
 954 => x"12",
 955 => x"F1",
 956 => x"AE",
 957 => x"C3",
 958 => x"AE",
 959 => x"EF",
 960 => x"90",
 961 => x"6F",
 962 => x"A2",
 963 => x"90",
 964 => x"6F",
 965 => x"C1",
 966 => x"16",
 967 => x"F1",
 968 => x"AE",
 969 => x"C3",
 970 => x"AE",
 971 => x"EF",
 972 => x"B0",
 973 => x"0B",
 974 => x"90",
 975 => x"61",
 976 => x"70",
 977 => x"72",
 978 => x"70",
 979 => x"90",
 980 => x"46",
 981 => x"61",
 982 => x"A6",
 983 => x"90",
 984 => x"60",
 985 => x"B0",
 986 => x"0E",
 987 => x"15",
 988 => x"16",
 989 => x"10",
 990 => x"15",
 991 => x"F1",
 992 => x"90",
 993 => x"61",
 994 => x"A6",
 995 => x"90",
 996 => x"71",
 997 => x"40",
 998 => x"61",
 999 => x"72",
1000 => x"9E",
1001 => x"61",
1002 => x"A6",
1003 => x"70",
1004 => x"06",
1005 => x"70",
1006 => x"36",
1007 => x"6F",
1008 => x"B0",
1009 => x"0B",
1010 => x"90",
1011 => x"61",
1012 => x"B0",
1013 => x"0E",
1014 => x"10",
1015 => x"F1",
1016 => x"90",
1017 => x"60",
1018 => x"90",
1019 => x"61",
1020 => x"B0",
1021 => x"0B",
1022 => x"90",
1023 => x"61",
1024 => x"70",
1025 => x"70",
1026 => x"90",
1027 => x"60",
1028 => x"34",
1029 => x"60",
1030 => x"A2",
1031 => x"70",
1032 => x"27",
1033 => x"30",
1034 => x"71",
1035 => x"71",
1036 => x"70",
1037 => x"40",
1038 => x"41",
1039 => x"00",
1040 => x"71",
1041 => x"40",
1042 => x"60",
1043 => x"B0",
1044 => x"0C",
1045 => x"90",
1046 => x"61",
1047 => x"72",
1048 => x"70",
1049 => x"90",
1050 => x"47",
1051 => x"61",
1052 => x"A7",
1053 => x"90",
1054 => x"60",
1055 => x"B0",
1056 => x"0E",
1057 => x"11",
1058 => x"17",
1059 => x"10",
1060 => x"11",
1061 => x"F1",
1062 => x"70",
1063 => x"90",
1064 => x"60",
1065 => x"34",
1066 => x"60",
1067 => x"E2",
1068 => x"F1",
1069 => x"AE",
1070 => x"C3",
1071 => x"AE",
1072 => x"EF",
1073 => x"90",
1074 => x"60",
1075 => x"73",
1076 => x"90",
1077 => x"61",
1078 => x"F1",
1079 => x"AE",
1080 => x"C3",
1081 => x"AE",
1082 => x"EF",
1083 => x"A3",
1084 => x"71",
1085 => x"24",
1086 => x"30",
1087 => x"60",
1088 => x"B0",
1089 => x"0B",
1090 => x"91",
1091 => x"60",
1092 => x"77",
1093 => x"90",
1094 => x"61",
1095 => x"73",
1096 => x"70",
1097 => x"90",
1098 => x"40",
1099 => x"61",
1100 => x"A4",
1101 => x"70",
1102 => x"40",
1103 => x"40",
1104 => x"00",
1105 => x"90",
1106 => x"60",
1107 => x"F1",
1108 => x"AE",
1109 => x"C3",
1110 => x"AE",
1111 => x"EF",
1112 => x"B0",
1113 => x"0C",
1114 => x"90",
1115 => x"60",
1116 => x"F1",
1117 => x"AE",
1118 => x"C3",
1119 => x"AE",
1120 => x"EF",
1121 => x"AE",
1122 => x"E5",
1123 => x"C0",
1124 => x"7F",
1125 => x"04",
1126 => x"90",
1127 => x"60",
1128 => x"A2",
1129 => x"7F",
1130 => x"05",
1131 => x"F1",
1132 => x"AE",
1133 => x"F1",
1134 => x"AE",
1135 => x"C0",
1136 => x"7F",
1137 => x"01",
1138 => x"24",
1139 => x"D0",
1140 => x"D0",
1141 => x"D0",
1142 => x"D0",
1143 => x"24",
1144 => x"C0",
1145 => x"C2",
1146 => x"02",
1147 => x"22",
1148 => x"72",
1149 => x"54",
1150 => x"22",
1151 => x"78",
1152 => x"54",
1153 => x"22",
1154 => x"B0",
1155 => x"FF",
1156 => x"02",
1157 => x"C3",
1158 => x"AE",
1159 => x"EF",
1160 => x"AE",
1161 => x"E9",
1162 => x"AE",
1163 => x"E8",
1164 => x"AE",
1165 => x"E7",
1166 => x"AE",
1167 => x"E6",
1168 => x"AE",
1169 => x"E5",
1170 => x"70",
1171 => x"A3",
1172 => x"70",
1173 => x"A4",
1174 => x"70",
1175 => x"70",
1176 => x"90",
1177 => x"60",
1178 => x"71",
1179 => x"22",
1180 => x"30",
1181 => x"60",
1182 => x"70",
1183 => x"22",
1184 => x"30",
1185 => x"60",
1186 => x"70",
1187 => x"22",
1188 => x"30",
1189 => x"60",
1190 => x"70",
1191 => x"22",
1192 => x"30",
1193 => x"60",
1194 => x"A2",
1195 => x"73",
1196 => x"40",
1197 => x"00",
1198 => x"70",
1199 => x"70",
1200 => x"40",
1201 => x"41",
1202 => x"00",
1203 => x"70",
1204 => x"C2",
1205 => x"32",
1206 => x"6F",
1207 => x"28",
1208 => x"30",
1209 => x"6F",
1210 => x"A7",
1211 => x"15",
1212 => x"15",
1213 => x"15",
1214 => x"15",
1215 => x"15",
1216 => x"9D",
1217 => x"60",
1218 => x"37",
1219 => x"6F",
1220 => x"D0",
1221 => x"D0",
1222 => x"D0",
1223 => x"D0",
1224 => x"A7",
1225 => x"B0",
1226 => x"0C",
1227 => x"9C",
1228 => x"60",
1229 => x"70",
1230 => x"60",
1231 => x"70",
1232 => x"A6",
1233 => x"37",
1234 => x"A6",
1235 => x"37",
1236 => x"60",
1237 => x"A7",
1238 => x"B0",
1239 => x"0C",
1240 => x"9F",
1241 => x"60",
1242 => x"34",
1243 => x"60",
1244 => x"A8",
1245 => x"A5",
1246 => x"90",
1247 => x"38",
1248 => x"60",
1249 => x"60",
1250 => x"38",
1251 => x"60",
1252 => x"60",
1253 => x"39",
1254 => x"6F",
1255 => x"A5",
1256 => x"F1",
1257 => x"AE",
1258 => x"F1",
1259 => x"AE",
1260 => x"F1",
1261 => x"AE",
1262 => x"F1",
1263 => x"AE",
1264 => x"F1",
1265 => x"AE",
1266 => x"F1",
1267 => x"AE",
1268 => x"C3",
1269 => x"AE",
1270 => x"EF",
1271 => x"C1",
1272 => x"90",
1273 => x"60",
1274 => x"C1",
1275 => x"F1",
1276 => x"AE",
1277 => x"AE",
1278 => x"EF",
1279 => x"C0",
1280 => x"90",
1281 => x"60",
1282 => x"C0",
1283 => x"F1",
1284 => x"AE",
1285 => x"D0",
1286 => x"D0",
1287 => x"D0",
1288 => x"D0",
1289 => x"70",
1290 => x"01",
1291 => x"73",
1292 => x"11",
1293 => x"73",
1294 => x"40",
1295 => x"A1",
1296 => x"F0",
1297 => x"30",
1298 => x"6F",
1299 => x"E1",
1300 => x"70",
1301 => x"03",
1302 => x"73",
1303 => x"11",
1304 => x"73",
1305 => x"40",
1306 => x"A1",
1307 => x"F0",
1308 => x"30",
1309 => x"6F",
1310 => x"E1",
1311 => x"C3",
1312 => x"AE",
1313 => x"EF",
1314 => x"90",
1315 => x"60",
1316 => x"A4",
1317 => x"90",
1318 => x"6F",
1319 => x"A5",
1320 => x"33",
1321 => x"60",
1322 => x"90",
1323 => x"60",
1324 => x"F1",
1325 => x"AE",
1326 => x"C3",
1327 => x"AE",
1328 => x"EF",
1329 => x"A3",
1330 => x"F3",
1331 => x"90",
1332 => x"60",
1333 => x"A2",
1334 => x"A4",
1335 => x"34",
1336 => x"6F",
1337 => x"F1",
1338 => x"AE",
1339 => x"C3",
1340 => x"AE",
1341 => x"EF",
1342 => x"AE",
1343 => x"E4",
1344 => x"13",
1345 => x"F3",
1346 => x"A2",
1347 => x"33",
1348 => x"60",
1349 => x"9F",
1350 => x"60",
1351 => x"F1",
1352 => x"AE",
1353 => x"F1",
1354 => x"AE",
1355 => x"C3",
1356 => x"70",
1357 => x"7F",
1358 => x"03",
1359 => x"70",
1360 => x"20",
1361 => x"30",
1362 => x"60",
1363 => x"F0",
1364 => x"30",
1365 => x"6F",
1366 => x"70",
1367 => x"E0",
1368 => x"F0",
1369 => x"30",
1370 => x"6F",
1371 => x"E3",
1372 => x"C3",
1373 => x"AE",
1374 => x"EF",
1375 => x"90",
1376 => x"60",
1377 => x"76",
1378 => x"42",
1379 => x"60",
1380 => x"72",
1381 => x"40",
1382 => x"00",
1383 => x"F1",
1384 => x"AE",
1385 => x"C3",
1386 => x"F0",
1387 => x"32",
1388 => x"6F",
1389 => x"AC",
1390 => x"E0",
1391 => x"7F",
1392 => x"02",
1393 => x"C3",
1394 => x"53",
1395 => x"65",
1396 => x"74",
1397 => x"32",
1398 => x"4D",
1399 => x"6E",
1400 => x"74",
1401 => x"72",
1402 => x"4C",
1403 => x"61",
1404 => x"65",
1405 => x"20",
1406 => x"30",
1407 => x"39",
1408 => x"2D",
1409 => x"65",
1410 => x"61",
1411 => x"00",
1412 => x"3E",
1413 => x"00",
1414 => x"0A",
1415 => x"20",
1416 => x"20",
1417 => x"20",
1418 => x"75",
1419 => x"70",
1420 => x"6D",
1421 => x"6D",
1422 => x"72",
1423 => x"0A",
1424 => x"4D",
1425 => x"2D",
1426 => x"4D",
1427 => x"64",
1428 => x"66",
1429 => x"20",
1430 => x"65",
1431 => x"6F",
1432 => x"79",
1433 => x"20",
1434 => x"20",
1435 => x"20",
1436 => x"6F",
1437 => x"28",
1438 => x"78",
1439 => x"63",
1440 => x"74",
1441 => x"29",
1442 => x"20",
1443 => x"20",
1444 => x"20",
1445 => x"65",
1446 => x"69",
1447 => x"74",
1448 => x"72",
1449 => x"0A",
1450 => x"42",
1451 => x"2D",
1452 => x"42",
1453 => x"75",
1454 => x"20",
1455 => x"61",
1456 => x"65",
1457 => x"73",
1458 => x"74",
1459 => x"20",
1460 => x"20",
1461 => x"20",
1462 => x"70",
1463 => x"6F",
1464 => x"64",
1465 => x"53",
1466 => x"45",
1467 => x"66",
1468 => x"6C",
1469 => x"20",
1470 => x"6F",
1471 => x"20",
1472 => x"65",
1473 => x"64",
1474 => x"61",
1475 => x"20",
1476 => x"72",
1477 => x"6D",
1478 => x"74",
1479 => x"0A",
1480 => x"44",
1481 => x"6D",
1482 => x"20",
1483 => x"42",
1484 => x"75",
1485 => x"0A",
1486 => x"47",
1487 => x"20",
1488 => x"4D",
1489 => x"64",
1490 => x"66",
1491 => x"20",
1492 => x"52",
1493 => x"67",
1494 => x"73",
1495 => x"65",
1496 => x"73",
1497 => x"00",
1498 => x"6F",
1499 => x"69",
1500 => x"79",
1501 => x"72",
1502 => x"67",
1503 => x"30",
1504 => x"31",
1505 => x"20",
1506 => x"43",
1507 => x"66",
1508 => x"72",
1509 => x"70",
1510 => x"29",
1511 => x"00",
1512 => x"69",
1513 => x"74",
1514 => x"00",
1515 => x"70",
1516 => x"6F",
1517 => x"64",
1518 => x"41",
1519 => x"61",
1520 => x"74",
1521 => x"6E",
1522 => x"20",
1523 => x"57",
1524 => x"2E",
1525 => x"2E",
1526 => x"20",
1527 => x"63",
1528 => x"00",
1529 => x"4C",
1530 => x"61",
1531 => x"65",
1532 => x"20",
1533 => x"20",
1534 => x"52",
1535 => x"3D",
1536 => x"0A",
1537 => x"55",
1538 => x"6C",
1539 => x"61",
1540 => x"20",
1541 => x"72",
1542 => x"6F",
1543 => x"20",
1544 => x"28",
1545 => x"20",
1546 => x"4B",
1547 => x"20",
1548 => x"52",
1549 => x"20",
1550 => x"41",
1551 => x"21",
1552 => x"53",
1553 => x"69",
1554 => x"63",
1555 => x"20",
1556 => x"6F",
1557 => x"6E",
1558 => x"77",
1559 => x"62",
1560 => x"75",
1561 => x"20",
1562 => x"61",
1563 => x"65",
1564 => x"20",
1565 => x"79",
1566 => x"65",
1567 => x"27",
1568 => x"27",
1569 => x"73",
1570 => x"76",
1571 => x"72",
1572 => x"6C",
1573 => x"74",
1574 => x"6D",
1575 => x"73",
1576 => x"74",
1577 => x"20",
1578 => x"65",
1579 => x"2E",
1580 => x"55",
1581 => x"52",
1582 => x"3D",
1583 => x"4E",
1584 => x"77",
1585 => x"55",
1586 => x"52",
1587 => x"20",
1588 => x"70",
1589 => x"65",
1590 => x"3D",
1591 => x"0A",
1592 => x"78",
1593 => x"63",
1594 => x"74",
1595 => x"20",
1596 => x"2E",
1597 => x"2E",
1598 => x"0A",
1599 => x"2C",
1600 => x"00",
1601 => x"20",
1602 => x"08",
1603 => x"08",
1604 => x"08",
1605 => x"20",
1606 => x"08",
1607 => x"00",
1608 => x"20",
1609 => x"20",
1610 => x"20",
1611 => x"20",
1612 => x"0A",
1613 => x"58",
1614 => x"72",
1615 => x"20",
1616 => x"61",
1617 => x"20",
1618 => x"65",
1619 => x"65",
1620 => x"20",
1621 => x"2D",
1622 => x"00",
1623 => x"FF",
1624 => x"00",
1625 => x"01",
1626 => x"6F",
1627 => x"20",
1628 => x"20",
1629 => x"F0",
1630 => x"00",
1631 => x"01",
1632 => x"6E",
1633 => x"20",
1634 => x"20",
1635 => x"F0",
1636 => x"10",
1637 => x"01",
1638 => x"64",
1639 => x"20",
1640 => x"20",
1641 => x"F0",
1642 => x"20",
1643 => x"01",
1644 => x"6F",
1645 => x"20",
1646 => x"20",
1647 => x"F0",
1648 => x"30",
1649 => x"01",
1650 => x"73",
1651 => x"73",
1652 => x"7A",
1653 => x"F0",
1654 => x"30",
1655 => x"01",
1656 => x"73",
1657 => x"73",
1658 => x"20",
1659 => x"F0",
1660 => x"30",
1661 => x"01",
1662 => x"69",
1663 => x"73",
1664 => x"7A",
1665 => x"F0",
1666 => x"30",
1667 => x"01",
1668 => x"69",
1669 => x"73",
1670 => x"20",
1671 => x"F0",
1672 => x"40",
1673 => x"01",
1674 => x"75",
1675 => x"73",
1676 => x"74",
1677 => x"F0",
1678 => x"50",
1679 => x"01",
1680 => x"75",
1681 => x"20",
1682 => x"20",
1683 => x"F0",
1684 => x"60",
1685 => x"01",
1686 => x"6A",
1687 => x"70",
1688 => x"20",
1689 => x"F0",
1690 => x"70",
1691 => x"01",
1692 => x"64",
1693 => x"20",
1694 => x"20",
1695 => x"F0",
1696 => x"80",
1697 => x"02",
1698 => x"6A",
1699 => x"70",
1700 => x"20",
1701 => x"F0",
1702 => x"90",
1703 => x"01",
1704 => x"65",
1705 => x"70",
1706 => x"20",
1707 => x"F0",
1708 => x"A0",
1709 => x"01",
1710 => x"6F",
1711 => x"20",
1712 => x"20",
1713 => x"F0",
1714 => x"A0",
1715 => x"01",
1716 => x"6E",
1717 => x"73",
1718 => x"20",
1719 => x"FF",
1720 => x"B0",
1721 => x"02",
1722 => x"64",
1723 => x"20",
1724 => x"20",
1725 => x"FF",
1726 => x"B1",
1727 => x"03",
1728 => x"64",
1729 => x"20",
1730 => x"20",
1731 => x"FF",
1732 => x"B2",
1733 => x"01",
1734 => x"65",
1735 => x"69",
1736 => x"20",
1737 => x"FF",
1738 => x"B3",
1739 => x"01",
1740 => x"65",
1741 => x"69",
1742 => x"20",
1743 => x"FF",
1744 => x"B4",
1745 => x"01",
1746 => x"65",
1747 => x"63",
1748 => x"20",
1749 => x"FF",
1750 => x"B5",
1751 => x"01",
1752 => x"65",
1753 => x"74",
1754 => x"20",
1755 => x"FF",
1756 => x"B6",
1757 => x"01",
1758 => x"65",
1759 => x"78",
1760 => x"20",
1761 => x"FF",
1762 => x"B7",
1763 => x"01",
1764 => x"65",
1765 => x"74",
1766 => x"20",
1767 => x"FF",
1768 => x"C0",
1769 => x"01",
1770 => x"77",
1771 => x"70",
1772 => x"20",
1773 => x"FF",
1774 => x"C1",
1775 => x"01",
1776 => x"77",
1777 => x"70",
1778 => x"20",
1779 => x"FF",
1780 => x"C2",
1781 => x"01",
1782 => x"6F",
1783 => x"20",
1784 => x"20",
1785 => x"FF",
1786 => x"C3",
1787 => x"01",
1788 => x"6A",
1789 => x"70",
1790 => x"20",
1791 => x"FF",
1792 => x"D0",
1793 => x"01",
1794 => x"73",
1795 => x"20",
1796 => x"20",
1797 => x"FF",
1798 => x"D1",
1799 => x"01",
1800 => x"73",
1801 => x"20",
1802 => x"20",
1803 => x"F0",
1804 => x"E0",
1805 => x"01",
1806 => x"6F",
1807 => x"77",
1808 => x"20",
1809 => x"F0",
1810 => x"E0",
1811 => x"01",
1812 => x"6F",
1813 => x"64",
1814 => x"20",
1815 => x"F0",
1816 => x"E0",
1817 => x"01",
1818 => x"6F",
1819 => x"62",
1820 => x"20",
1821 => x"FF",
1822 => x"F0",
1823 => x"01",
1824 => x"6F",
1825 => x"77",
1826 => x"20",
1827 => x"FF",
1828 => x"F1",
1829 => x"01",
1830 => x"6F",
1831 => x"64",
1832 => x"20",
1833 => x"FF",
1834 => x"F2",
1835 => x"01",
1836 => x"6F",
1837 => x"73",
1838 => x"20",
1839 => x"FF",
1840 => x"F3",
1841 => x"01",
1842 => x"6F",
1843 => x"62",
1844 => x"20",
1845 => x"00",
1846 => x"00",
1847 => x"01",
1848 => x"3F",
1849 => x"20",
1850 => x"20",
1851 => x"30",
1852 => x"00",
1853 => x"00",
1854 => x"00",
1855 => x"00",
1856 => x"00",
1857 => x"00",
1858 => x"00",
1859 => x"00",
1860 => x"00",
1861 => x"00",
1862 => x"00",
1863 => x"00",
1864 => x"00",
1865 => x"00",
1866 => x"00",
1867 => x"00",
1868 => x"00",
1869 => x"00",
1870 => x"00",
1871 => x"00",
1872 => x"00",
1873 => x"00",
1874 => x"00",
1875 => x"00",
1876 => x"00",
1877 => x"00",
1878 => x"00",
1879 => x"00",
1880 => x"00",
1881 => x"00",
1882 => x"00",
1883 => x"00",
1884 => x"00",
1885 => x"00",
1886 => x"00",
1887 => x"00",
1888 => x"00",
1889 => x"00",
1890 => x"00",
1891 => x"00",
1892 => x"00",
1893 => x"00",
1894 => x"00",
1895 => x"00",
1896 => x"00",
1897 => x"00",
1898 => x"00",
1899 => x"00",
1900 => x"00",
1901 => x"00",
1902 => x"00",
1903 => x"00",
1904 => x"00",
1905 => x"00",
1906 => x"00",
1907 => x"00",
1908 => x"00",
1909 => x"00",
1910 => x"00",
1911 => x"00",
1912 => x"00",
1913 => x"00",
1914 => x"00",
1915 => x"00",
1916 => x"00",
1917 => x"00",
1918 => x"00",
1919 => x"00",
1920 => x"00",
1921 => x"00",
1922 => x"00",
1923 => x"00",
1924 => x"00",
1925 => x"00",
1926 => x"00",
1927 => x"00",
1928 => x"00",
1929 => x"00",
1930 => x"00",
1931 => x"00",
1932 => x"00",
1933 => x"00",
1934 => x"00",
1935 => x"00",
1936 => x"00",
1937 => x"00",
1938 => x"00",
1939 => x"00",
1940 => x"00",
1941 => x"00",
1942 => x"00",
1943 => x"00",
1944 => x"00",
1945 => x"00",
1946 => x"00",
1947 => x"00",
1948 => x"00",
1949 => x"00",
1950 => x"BA",
1951 => x"C0",


others => x"00"
);

attribute syn_ramstyle : string;
attribute syn_ramstyle of RAM : signal is "block_ram";

begin
   --busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(conv_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(conv_integer(addr_r));
end architecture behavioral; -- Entity: Sweet32_ROM