-- from http://help.latticesemi.com/docs/webhelp/eng/wwhelp/wwhimpl/common/html/wwhelp.htm#href=Design%20Entry/inferring_ram_dual_port.htm
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
 
entity font_dp_ram is
generic (
	addr_width : natural;
	data_width : natural);
port (
	addra_i	: in std_logic_vector (addr_width - 1 downto 0);
	wea_i	: in std_logic;
	clka_i	: in std_logic;
	dina_i	: in std_logic_vector (data_width - 1 downto 0);
	douta_o	: out std_logic_vector (data_width - 1 downto 0);
	addrb_i	: in std_logic_vector (addr_width - 1 downto 0);
	web_i	: in std_logic;
	clkb_i	: in std_logic;
	dinb_i	: in std_logic_vector (data_width - 1 downto 0);
	doutb_o	: out std_logic_vector (data_width - 1 downto 0));
end font_dp_ram;
 
architecture rtl of font_dp_ram is
	type mem_type is array ((2** addr_width) - 1 downto 0) of 
	std_logic_vector(data_width - 1 downto 0);
	signal mem : mem_type := (
   0 => x"7E",
   1 => x"C3",
   2 => x"99",
   3 => x"99",
   4 => x"F3",
   5 => x"E7",
   6 => x"E7",
   7 => x"FF",
   8 => x"E7",
   9 => x"E7",
  10 => x"7E",
  11 => x"00",
  12 => x"00",
  13 => x"00",
  14 => x"00",
  15 => x"76",
  16 => x"DC",
  17 => x"00",
  18 => x"76",
  19 => x"DC",
  20 => x"00",
  21 => x"00",
  22 => x"00",
  23 => x"00",
  24 => x"6E",
  25 => x"D8",
  26 => x"D8",
  27 => x"D8",
  28 => x"D8",
  29 => x"DE",
  30 => x"D8",
  31 => x"D8",
  32 => x"D8",
  33 => x"6E",
  34 => x"00",
  35 => x"00",
  36 => x"00",
  37 => x"00",
  38 => x"00",
  39 => x"6E",
  40 => x"DB",
  41 => x"DB",
  42 => x"DF",
  43 => x"D8",
  44 => x"DB",
  45 => x"6E",
  46 => x"00",
  47 => x"00",
  48 => x"00",
  49 => x"00",
  50 => x"10",
  51 => x"38",
  52 => x"7C",
  53 => x"FE",
  54 => x"7C",
  55 => x"38",
  56 => x"10",
  57 => x"00",
  58 => x"00",
  59 => x"00",
  60 => x"88",
  61 => x"88",
  62 => x"F8",
  63 => x"88",
  64 => x"88",
  65 => x"00",
  66 => x"3E",
  67 => x"08",
  68 => x"08",
  69 => x"08",
  70 => x"08",
  71 => x"00",
  72 => x"F8",
  73 => x"80",
  74 => x"E0",
  75 => x"80",
  76 => x"80",
  77 => x"00",
  78 => x"3E",
  79 => x"20",
  80 => x"38",
  81 => x"20",
  82 => x"20",
  83 => x"00",
  84 => x"78",
  85 => x"80",
  86 => x"80",
  87 => x"80",
  88 => x"78",
  89 => x"00",
  90 => x"3C",
  91 => x"22",
  92 => x"3E",
  93 => x"24",
  94 => x"22",
  95 => x"00",
  96 => x"80",
  97 => x"80",
  98 => x"80",
  99 => x"80",
 100 => x"F8",
 101 => x"00",
 102 => x"3E",
 103 => x"20",
 104 => x"38",
 105 => x"20",
 106 => x"20",
 107 => x"00",
 108 => x"22",
 109 => x"88",
 110 => x"22",
 111 => x"88",
 112 => x"22",
 113 => x"88",
 114 => x"22",
 115 => x"88",
 116 => x"22",
 117 => x"88",
 118 => x"22",
 119 => x"88",
 120 => x"55",
 121 => x"AA",
 122 => x"55",
 123 => x"AA",
 124 => x"55",
 125 => x"AA",
 126 => x"55",
 127 => x"AA",
 128 => x"55",
 129 => x"AA",
 130 => x"55",
 131 => x"AA",
 132 => x"EE",
 133 => x"BB",
 134 => x"EE",
 135 => x"BB",
 136 => x"EE",
 137 => x"BB",
 138 => x"EE",
 139 => x"BB",
 140 => x"EE",
 141 => x"BB",
 142 => x"EE",
 143 => x"BB",
 144 => x"FF",
 145 => x"FF",
 146 => x"FF",
 147 => x"FF",
 148 => x"FF",
 149 => x"FF",
 150 => x"FF",
 151 => x"FF",
 152 => x"FF",
 153 => x"FF",
 154 => x"FF",
 155 => x"FF",
 156 => x"00",
 157 => x"00",
 158 => x"00",
 159 => x"00",
 160 => x"00",
 161 => x"00",
 162 => x"FF",
 163 => x"FF",
 164 => x"FF",
 165 => x"FF",
 166 => x"FF",
 167 => x"FF",
 168 => x"FF",
 169 => x"FF",
 170 => x"FF",
 171 => x"FF",
 172 => x"FF",
 173 => x"FF",
 174 => x"00",
 175 => x"00",
 176 => x"00",
 177 => x"00",
 178 => x"00",
 179 => x"00",
 180 => x"F0",
 181 => x"F0",
 182 => x"F0",
 183 => x"F0",
 184 => x"F0",
 185 => x"F0",
 186 => x"F0",
 187 => x"F0",
 188 => x"F0",
 189 => x"F0",
 190 => x"F0",
 191 => x"F0",
 192 => x"0F",
 193 => x"0F",
 194 => x"0F",
 195 => x"0F",
 196 => x"0F",
 197 => x"0F",
 198 => x"0F",
 199 => x"0F",
 200 => x"0F",
 201 => x"0F",
 202 => x"0F",
 203 => x"0F",
 204 => x"88",
 205 => x"C8",
 206 => x"A8",
 207 => x"98",
 208 => x"88",
 209 => x"00",
 210 => x"20",
 211 => x"20",
 212 => x"20",
 213 => x"20",
 214 => x"3E",
 215 => x"00",
 216 => x"88",
 217 => x"88",
 218 => x"50",
 219 => x"50",
 220 => x"20",
 221 => x"00",
 222 => x"3E",
 223 => x"08",
 224 => x"08",
 225 => x"08",
 226 => x"08",
 227 => x"00",
 228 => x"00",
 229 => x"00",
 230 => x"06",
 231 => x"0C",
 232 => x"18",
 233 => x"30",
 234 => x"7E",
 235 => x"00",
 236 => x"7E",
 237 => x"00",
 238 => x"00",
 239 => x"00",
 240 => x"00",
 241 => x"00",
 242 => x"60",
 243 => x"30",
 244 => x"18",
 245 => x"0C",
 246 => x"7E",
 247 => x"00",
 248 => x"7E",
 249 => x"00",
 250 => x"00",
 251 => x"00",
 252 => x"00",
 253 => x"00",
 254 => x"06",
 255 => x"0C",
 256 => x"FE",
 257 => x"38",
 258 => x"FE",
 259 => x"60",
 260 => x"C0",
 261 => x"00",
 262 => x"00",
 263 => x"00",
 264 => x"00",
 265 => x"02",
 266 => x"0E",
 267 => x"3E",
 268 => x"7E",
 269 => x"FE",
 270 => x"7E",
 271 => x"3E",
 272 => x"0E",
 273 => x"02",
 274 => x"00",
 275 => x"00",
 276 => x"00",
 277 => x"80",
 278 => x"E0",
 279 => x"F0",
 280 => x"FC",
 281 => x"FE",
 282 => x"FC",
 283 => x"F0",
 284 => x"E0",
 285 => x"80",
 286 => x"00",
 287 => x"00",
 288 => x"00",
 289 => x"18",
 290 => x"3C",
 291 => x"7E",
 292 => x"18",
 293 => x"18",
 294 => x"18",
 295 => x"18",
 296 => x"18",
 297 => x"18",
 298 => x"00",
 299 => x"00",
 300 => x"00",
 301 => x"18",
 302 => x"18",
 303 => x"18",
 304 => x"18",
 305 => x"18",
 306 => x"18",
 307 => x"7E",
 308 => x"3C",
 309 => x"18",
 310 => x"00",
 311 => x"00",
 312 => x"00",
 313 => x"00",
 314 => x"00",
 315 => x"18",
 316 => x"0C",
 317 => x"FE",
 318 => x"0C",
 319 => x"18",
 320 => x"00",
 321 => x"00",
 322 => x"00",
 323 => x"00",
 324 => x"00",
 325 => x"00",
 326 => x"00",
 327 => x"30",
 328 => x"60",
 329 => x"FE",
 330 => x"60",
 331 => x"30",
 332 => x"00",
 333 => x"00",
 334 => x"00",
 335 => x"00",
 336 => x"00",
 337 => x"18",
 338 => x"3C",
 339 => x"7E",
 340 => x"18",
 341 => x"18",
 342 => x"18",
 343 => x"7E",
 344 => x"3C",
 345 => x"18",
 346 => x"00",
 347 => x"00",
 348 => x"00",
 349 => x"00",
 350 => x"00",
 351 => x"28",
 352 => x"6C",
 353 => x"FE",
 354 => x"6C",
 355 => x"28",
 356 => x"00",
 357 => x"00",
 358 => x"00",
 359 => x"00",
 360 => x"00",
 361 => x"06",
 362 => x"06",
 363 => x"36",
 364 => x"66",
 365 => x"FE",
 366 => x"60",
 367 => x"30",
 368 => x"00",
 369 => x"00",
 370 => x"00",
 371 => x"00",
 372 => x"00",
 373 => x"00",
 374 => x"00",
 375 => x"C0",
 376 => x"7C",
 377 => x"6E",
 378 => x"6C",
 379 => x"6C",
 380 => x"6C",
 381 => x"00",
 382 => x"00",
 383 => x"00",
 384 => x"00",
 385 => x"00",
 386 => x"00",
 387 => x"00",
 388 => x"00",
 389 => x"00",
 390 => x"00",
 391 => x"00",
 392 => x"00",
 393 => x"00",
 394 => x"00",
 395 => x"00",
 396 => x"00",
 397 => x"18",
 398 => x"3C",
 399 => x"3C",
 400 => x"3C",
 401 => x"18",
 402 => x"18",
 403 => x"00",
 404 => x"18",
 405 => x"18",
 406 => x"00",
 407 => x"00",
 408 => x"00",
 409 => x"36",
 410 => x"36",
 411 => x"14",
 412 => x"00",
 413 => x"00",
 414 => x"00",
 415 => x"00",
 416 => x"00",
 417 => x"00",
 418 => x"00",
 419 => x"00",
 420 => x"00",
 421 => x"00",
 422 => x"00",
 423 => x"6C",
 424 => x"FE",
 425 => x"6C",
 426 => x"6C",
 427 => x"6C",
 428 => x"FE",
 429 => x"6C",
 430 => x"00",
 431 => x"00",
 432 => x"00",
 433 => x"10",
 434 => x"7C",
 435 => x"D6",
 436 => x"70",
 437 => x"38",
 438 => x"1C",
 439 => x"D6",
 440 => x"7C",
 441 => x"10",
 442 => x"00",
 443 => x"00",
 444 => x"00",
 445 => x"00",
 446 => x"00",
 447 => x"62",
 448 => x"66",
 449 => x"0C",
 450 => x"18",
 451 => x"30",
 452 => x"66",
 453 => x"C6",
 454 => x"00",
 455 => x"00",
 456 => x"00",
 457 => x"38",
 458 => x"6C",
 459 => x"38",
 460 => x"38",
 461 => x"72",
 462 => x"FE",
 463 => x"CC",
 464 => x"CC",
 465 => x"76",
 466 => x"00",
 467 => x"00",
 468 => x"1C",
 469 => x"1C",
 470 => x"0C",
 471 => x"18",
 472 => x"00",
 473 => x"00",
 474 => x"00",
 475 => x"00",
 476 => x"00",
 477 => x"00",
 478 => x"00",
 479 => x"00",
 480 => x"00",
 481 => x"0C",
 482 => x"18",
 483 => x"30",
 484 => x"30",
 485 => x"30",
 486 => x"30",
 487 => x"30",
 488 => x"18",
 489 => x"0C",
 490 => x"00",
 491 => x"00",
 492 => x"00",
 493 => x"30",
 494 => x"18",
 495 => x"0C",
 496 => x"0C",
 497 => x"0C",
 498 => x"0C",
 499 => x"0C",
 500 => x"18",
 501 => x"30",
 502 => x"00",
 503 => x"00",
 504 => x"00",
 505 => x"00",
 506 => x"00",
 507 => x"6C",
 508 => x"38",
 509 => x"FE",
 510 => x"38",
 511 => x"6C",
 512 => x"00",
 513 => x"00",
 514 => x"00",
 515 => x"00",
 516 => x"00",
 517 => x"00",
 518 => x"00",
 519 => x"18",
 520 => x"18",
 521 => x"7E",
 522 => x"18",
 523 => x"18",
 524 => x"00",
 525 => x"00",
 526 => x"00",
 527 => x"00",
 528 => x"00",
 529 => x"00",
 530 => x"00",
 531 => x"00",
 532 => x"00",
 533 => x"00",
 534 => x"00",
 535 => x"0C",
 536 => x"0C",
 537 => x"0C",
 538 => x"18",
 539 => x"00",
 540 => x"00",
 541 => x"00",
 542 => x"00",
 543 => x"00",
 544 => x"00",
 545 => x"FE",
 546 => x"00",
 547 => x"00",
 548 => x"00",
 549 => x"00",
 550 => x"00",
 551 => x"00",
 552 => x"00",
 553 => x"00",
 554 => x"00",
 555 => x"00",
 556 => x"00",
 557 => x"00",
 558 => x"00",
 559 => x"00",
 560 => x"18",
 561 => x"18",
 562 => x"00",
 563 => x"00",
 564 => x"00",
 565 => x"00",
 566 => x"00",
 567 => x"06",
 568 => x"0C",
 569 => x"18",
 570 => x"30",
 571 => x"60",
 572 => x"C0",
 573 => x"00",
 574 => x"00",
 575 => x"00",
 576 => x"00",
 577 => x"7C",
 578 => x"C6",
 579 => x"C6",
 580 => x"C6",
 581 => x"D6",
 582 => x"C6",
 583 => x"C6",
 584 => x"C6",
 585 => x"7C",
 586 => x"00",
 587 => x"00",
 588 => x"00",
 589 => x"18",
 590 => x"78",
 591 => x"18",
 592 => x"18",
 593 => x"18",
 594 => x"18",
 595 => x"18",
 596 => x"18",
 597 => x"7E",
 598 => x"00",
 599 => x"00",
 600 => x"00",
 601 => x"7C",
 602 => x"C6",
 603 => x"C6",
 604 => x"0C",
 605 => x"18",
 606 => x"30",
 607 => x"60",
 608 => x"C6",
 609 => x"FE",
 610 => x"00",
 611 => x"00",
 612 => x"00",
 613 => x"7C",
 614 => x"C6",
 615 => x"06",
 616 => x"06",
 617 => x"3C",
 618 => x"06",
 619 => x"06",
 620 => x"C6",
 621 => x"7C",
 622 => x"00",
 623 => x"00",
 624 => x"00",
 625 => x"0C",
 626 => x"1C",
 627 => x"3C",
 628 => x"6C",
 629 => x"CC",
 630 => x"FE",
 631 => x"0C",
 632 => x"0C",
 633 => x"0C",
 634 => x"00",
 635 => x"00",
 636 => x"00",
 637 => x"FE",
 638 => x"C0",
 639 => x"C0",
 640 => x"C0",
 641 => x"FC",
 642 => x"06",
 643 => x"06",
 644 => x"C6",
 645 => x"7C",
 646 => x"00",
 647 => x"00",
 648 => x"00",
 649 => x"7C",
 650 => x"C6",
 651 => x"C0",
 652 => x"C0",
 653 => x"FC",
 654 => x"C6",
 655 => x"C6",
 656 => x"C6",
 657 => x"7C",
 658 => x"00",
 659 => x"00",
 660 => x"00",
 661 => x"FE",
 662 => x"C6",
 663 => x"0C",
 664 => x"18",
 665 => x"30",
 666 => x"30",
 667 => x"30",
 668 => x"30",
 669 => x"30",
 670 => x"00",
 671 => x"00",
 672 => x"00",
 673 => x"7C",
 674 => x"C6",
 675 => x"C6",
 676 => x"C6",
 677 => x"7C",
 678 => x"C6",
 679 => x"C6",
 680 => x"C6",
 681 => x"7C",
 682 => x"00",
 683 => x"00",
 684 => x"00",
 685 => x"7C",
 686 => x"C6",
 687 => x"C6",
 688 => x"C6",
 689 => x"7E",
 690 => x"06",
 691 => x"06",
 692 => x"C6",
 693 => x"7C",
 694 => x"00",
 695 => x"00",
 696 => x"00",
 697 => x"00",
 698 => x"00",
 699 => x"0C",
 700 => x"0C",
 701 => x"00",
 702 => x"00",
 703 => x"0C",
 704 => x"0C",
 705 => x"00",
 706 => x"00",
 707 => x"00",
 708 => x"00",
 709 => x"00",
 710 => x"00",
 711 => x"0C",
 712 => x"0C",
 713 => x"00",
 714 => x"00",
 715 => x"0C",
 716 => x"0C",
 717 => x"0C",
 718 => x"18",
 719 => x"00",
 720 => x"00",
 721 => x"0C",
 722 => x"18",
 723 => x"30",
 724 => x"60",
 725 => x"C0",
 726 => x"60",
 727 => x"30",
 728 => x"18",
 729 => x"0C",
 730 => x"00",
 731 => x"00",
 732 => x"00",
 733 => x"00",
 734 => x"00",
 735 => x"00",
 736 => x"FE",
 737 => x"00",
 738 => x"FE",
 739 => x"00",
 740 => x"00",
 741 => x"00",
 742 => x"00",
 743 => x"00",
 744 => x"00",
 745 => x"60",
 746 => x"30",
 747 => x"18",
 748 => x"0C",
 749 => x"06",
 750 => x"0C",
 751 => x"18",
 752 => x"30",
 753 => x"60",
 754 => x"00",
 755 => x"00",
 756 => x"00",
 757 => x"7C",
 758 => x"C6",
 759 => x"C6",
 760 => x"0C",
 761 => x"18",
 762 => x"18",
 763 => x"00",
 764 => x"18",
 765 => x"18",
 766 => x"00",
 767 => x"00",
 768 => x"00",
 769 => x"7C",
 770 => x"C6",
 771 => x"C6",
 772 => x"DE",
 773 => x"DE",
 774 => x"DE",
 775 => x"DC",
 776 => x"C0",
 777 => x"7E",
 778 => x"00",
 779 => x"00",
 780 => x"00",
 781 => x"38",
 782 => x"6C",
 783 => x"C6",
 784 => x"C6",
 785 => x"C6",
 786 => x"FE",
 787 => x"C6",
 788 => x"C6",
 789 => x"C6",
 790 => x"00",
 791 => x"00",
 792 => x"00",
 793 => x"FC",
 794 => x"66",
 795 => x"66",
 796 => x"66",
 797 => x"7C",
 798 => x"66",
 799 => x"66",
 800 => x"66",
 801 => x"FC",
 802 => x"00",
 803 => x"00",
 804 => x"00",
 805 => x"3C",
 806 => x"66",
 807 => x"C0",
 808 => x"C0",
 809 => x"C0",
 810 => x"C0",
 811 => x"C0",
 812 => x"66",
 813 => x"3C",
 814 => x"00",
 815 => x"00",
 816 => x"00",
 817 => x"F8",
 818 => x"6C",
 819 => x"66",
 820 => x"66",
 821 => x"66",
 822 => x"66",
 823 => x"66",
 824 => x"6C",
 825 => x"F8",
 826 => x"00",
 827 => x"00",
 828 => x"00",
 829 => x"FE",
 830 => x"66",
 831 => x"60",
 832 => x"60",
 833 => x"7C",
 834 => x"60",
 835 => x"60",
 836 => x"66",
 837 => x"FE",
 838 => x"00",
 839 => x"00",
 840 => x"00",
 841 => x"FE",
 842 => x"66",
 843 => x"60",
 844 => x"60",
 845 => x"7C",
 846 => x"60",
 847 => x"60",
 848 => x"60",
 849 => x"F0",
 850 => x"00",
 851 => x"00",
 852 => x"00",
 853 => x"7C",
 854 => x"C6",
 855 => x"C6",
 856 => x"C0",
 857 => x"C0",
 858 => x"CE",
 859 => x"C6",
 860 => x"C6",
 861 => x"7C",
 862 => x"00",
 863 => x"00",
 864 => x"00",
 865 => x"C6",
 866 => x"C6",
 867 => x"C6",
 868 => x"C6",
 869 => x"FE",
 870 => x"C6",
 871 => x"C6",
 872 => x"C6",
 873 => x"C6",
 874 => x"00",
 875 => x"00",
 876 => x"00",
 877 => x"3C",
 878 => x"18",
 879 => x"18",
 880 => x"18",
 881 => x"18",
 882 => x"18",
 883 => x"18",
 884 => x"18",
 885 => x"3C",
 886 => x"00",
 887 => x"00",
 888 => x"00",
 889 => x"3C",
 890 => x"18",
 891 => x"18",
 892 => x"18",
 893 => x"18",
 894 => x"18",
 895 => x"D8",
 896 => x"D8",
 897 => x"70",
 898 => x"00",
 899 => x"00",
 900 => x"00",
 901 => x"C6",
 902 => x"CC",
 903 => x"D8",
 904 => x"F0",
 905 => x"F0",
 906 => x"D8",
 907 => x"CC",
 908 => x"C6",
 909 => x"C6",
 910 => x"00",
 911 => x"00",
 912 => x"00",
 913 => x"F0",
 914 => x"60",
 915 => x"60",
 916 => x"60",
 917 => x"60",
 918 => x"60",
 919 => x"62",
 920 => x"66",
 921 => x"FE",
 922 => x"00",
 923 => x"00",
 924 => x"00",
 925 => x"C6",
 926 => x"C6",
 927 => x"EE",
 928 => x"FE",
 929 => x"D6",
 930 => x"D6",
 931 => x"D6",
 932 => x"C6",
 933 => x"C6",
 934 => x"00",
 935 => x"00",
 936 => x"00",
 937 => x"C6",
 938 => x"C6",
 939 => x"E6",
 940 => x"E6",
 941 => x"F6",
 942 => x"DE",
 943 => x"CE",
 944 => x"CE",
 945 => x"C6",
 946 => x"00",
 947 => x"00",
 948 => x"00",
 949 => x"7C",
 950 => x"C6",
 951 => x"C6",
 952 => x"C6",
 953 => x"C6",
 954 => x"C6",
 955 => x"C6",
 956 => x"C6",
 957 => x"7C",
 958 => x"00",
 959 => x"00",
 960 => x"00",
 961 => x"FC",
 962 => x"66",
 963 => x"66",
 964 => x"66",
 965 => x"7C",
 966 => x"60",
 967 => x"60",
 968 => x"60",
 969 => x"F0",
 970 => x"00",
 971 => x"00",
 972 => x"00",
 973 => x"7C",
 974 => x"C6",
 975 => x"C6",
 976 => x"C6",
 977 => x"C6",
 978 => x"C6",
 979 => x"C6",
 980 => x"D6",
 981 => x"7C",
 982 => x"06",
 983 => x"00",
 984 => x"00",
 985 => x"FC",
 986 => x"66",
 987 => x"66",
 988 => x"66",
 989 => x"7C",
 990 => x"78",
 991 => x"6C",
 992 => x"66",
 993 => x"E6",
 994 => x"00",
 995 => x"00",
 996 => x"00",
 997 => x"7C",
 998 => x"C6",
 999 => x"C0",
1000 => x"60",
1001 => x"38",
1002 => x"0C",
1003 => x"06",
1004 => x"C6",
1005 => x"7C",
1006 => x"00",
1007 => x"00",
1008 => x"00",
1009 => x"7E",
1010 => x"5A",
1011 => x"18",
1012 => x"18",
1013 => x"18",
1014 => x"18",
1015 => x"18",
1016 => x"18",
1017 => x"3C",
1018 => x"00",
1019 => x"00",
1020 => x"00",
1021 => x"C6",
1022 => x"C6",
1023 => x"C6",
1024 => x"C6",
1025 => x"C6",
1026 => x"C6",
1027 => x"C6",
1028 => x"C6",
1029 => x"7C",
1030 => x"00",
1031 => x"00",
1032 => x"00",
1033 => x"C6",
1034 => x"C6",
1035 => x"C6",
1036 => x"C6",
1037 => x"C6",
1038 => x"C6",
1039 => x"6C",
1040 => x"38",
1041 => x"10",
1042 => x"00",
1043 => x"00",
1044 => x"00",
1045 => x"C6",
1046 => x"C6",
1047 => x"D6",
1048 => x"D6",
1049 => x"D6",
1050 => x"FE",
1051 => x"EE",
1052 => x"C6",
1053 => x"C6",
1054 => x"00",
1055 => x"00",
1056 => x"00",
1057 => x"C6",
1058 => x"C6",
1059 => x"6C",
1060 => x"38",
1061 => x"38",
1062 => x"38",
1063 => x"6C",
1064 => x"C6",
1065 => x"C6",
1066 => x"00",
1067 => x"00",
1068 => x"00",
1069 => x"66",
1070 => x"66",
1071 => x"66",
1072 => x"66",
1073 => x"3C",
1074 => x"18",
1075 => x"18",
1076 => x"18",
1077 => x"3C",
1078 => x"00",
1079 => x"00",
1080 => x"00",
1081 => x"FE",
1082 => x"C6",
1083 => x"8C",
1084 => x"18",
1085 => x"30",
1086 => x"60",
1087 => x"C2",
1088 => x"C6",
1089 => x"FE",
1090 => x"00",
1091 => x"00",
1092 => x"00",
1093 => x"7C",
1094 => x"60",
1095 => x"60",
1096 => x"60",
1097 => x"60",
1098 => x"60",
1099 => x"60",
1100 => x"60",
1101 => x"7C",
1102 => x"00",
1103 => x"00",
1104 => x"00",
1105 => x"00",
1106 => x"00",
1107 => x"C0",
1108 => x"60",
1109 => x"30",
1110 => x"18",
1111 => x"0C",
1112 => x"06",
1113 => x"00",
1114 => x"00",
1115 => x"00",
1116 => x"00",
1117 => x"7C",
1118 => x"0C",
1119 => x"0C",
1120 => x"0C",
1121 => x"0C",
1122 => x"0C",
1123 => x"0C",
1124 => x"0C",
1125 => x"7C",
1126 => x"00",
1127 => x"00",
1128 => x"00",
1129 => x"18",
1130 => x"3C",
1131 => x"66",
1132 => x"00",
1133 => x"00",
1134 => x"00",
1135 => x"00",
1136 => x"00",
1137 => x"00",
1138 => x"00",
1139 => x"00",
1140 => x"00",
1141 => x"00",
1142 => x"00",
1143 => x"00",
1144 => x"00",
1145 => x"00",
1146 => x"00",
1147 => x"00",
1148 => x"00",
1149 => x"00",
1150 => x"00",
1151 => x"FF",
1152 => x"1C",
1153 => x"1C",
1154 => x"18",
1155 => x"0C",
1156 => x"00",
1157 => x"00",
1158 => x"00",
1159 => x"00",
1160 => x"00",
1161 => x"00",
1162 => x"00",
1163 => x"00",
1164 => x"00",
1165 => x"00",
1166 => x"00",
1167 => x"00",
1168 => x"78",
1169 => x"0C",
1170 => x"7C",
1171 => x"CC",
1172 => x"DC",
1173 => x"76",
1174 => x"00",
1175 => x"00",
1176 => x"00",
1177 => x"E0",
1178 => x"60",
1179 => x"60",
1180 => x"7C",
1181 => x"66",
1182 => x"66",
1183 => x"66",
1184 => x"66",
1185 => x"FC",
1186 => x"00",
1187 => x"00",
1188 => x"00",
1189 => x"00",
1190 => x"00",
1191 => x"00",
1192 => x"7C",
1193 => x"C6",
1194 => x"C0",
1195 => x"C0",
1196 => x"C6",
1197 => x"7C",
1198 => x"00",
1199 => x"00",
1200 => x"00",
1201 => x"1C",
1202 => x"0C",
1203 => x"0C",
1204 => x"7C",
1205 => x"CC",
1206 => x"CC",
1207 => x"CC",
1208 => x"CC",
1209 => x"7E",
1210 => x"00",
1211 => x"00",
1212 => x"00",
1213 => x"00",
1214 => x"00",
1215 => x"00",
1216 => x"7C",
1217 => x"C6",
1218 => x"FE",
1219 => x"C0",
1220 => x"C6",
1221 => x"7C",
1222 => x"00",
1223 => x"00",
1224 => x"00",
1225 => x"1C",
1226 => x"36",
1227 => x"30",
1228 => x"30",
1229 => x"FC",
1230 => x"30",
1231 => x"30",
1232 => x"30",
1233 => x"78",
1234 => x"00",
1235 => x"00",
1236 => x"00",
1237 => x"00",
1238 => x"00",
1239 => x"00",
1240 => x"76",
1241 => x"CE",
1242 => x"C6",
1243 => x"C6",
1244 => x"7E",
1245 => x"06",
1246 => x"C6",
1247 => x"7C",
1248 => x"00",
1249 => x"E0",
1250 => x"60",
1251 => x"60",
1252 => x"6C",
1253 => x"76",
1254 => x"66",
1255 => x"66",
1256 => x"66",
1257 => x"E6",
1258 => x"00",
1259 => x"00",
1260 => x"00",
1261 => x"18",
1262 => x"18",
1263 => x"00",
1264 => x"38",
1265 => x"18",
1266 => x"18",
1267 => x"18",
1268 => x"18",
1269 => x"3C",
1270 => x"00",
1271 => x"00",
1272 => x"00",
1273 => x"00",
1274 => x"0C",
1275 => x"0C",
1276 => x"00",
1277 => x"1C",
1278 => x"0C",
1279 => x"0C",
1280 => x"0C",
1281 => x"CC",
1282 => x"CC",
1283 => x"78",
1284 => x"00",
1285 => x"E0",
1286 => x"60",
1287 => x"60",
1288 => x"66",
1289 => x"6C",
1290 => x"78",
1291 => x"6C",
1292 => x"66",
1293 => x"E6",
1294 => x"00",
1295 => x"00",
1296 => x"00",
1297 => x"70",
1298 => x"30",
1299 => x"30",
1300 => x"30",
1301 => x"30",
1302 => x"30",
1303 => x"30",
1304 => x"34",
1305 => x"18",
1306 => x"00",
1307 => x"00",
1308 => x"00",
1309 => x"00",
1310 => x"00",
1311 => x"00",
1312 => x"6C",
1313 => x"FE",
1314 => x"D6",
1315 => x"D6",
1316 => x"C6",
1317 => x"C6",
1318 => x"00",
1319 => x"00",
1320 => x"00",
1321 => x"00",
1322 => x"00",
1323 => x"00",
1324 => x"DC",
1325 => x"66",
1326 => x"66",
1327 => x"66",
1328 => x"66",
1329 => x"66",
1330 => x"00",
1331 => x"00",
1332 => x"00",
1333 => x"00",
1334 => x"00",
1335 => x"00",
1336 => x"7C",
1337 => x"C6",
1338 => x"C6",
1339 => x"C6",
1340 => x"C6",
1341 => x"7C",
1342 => x"00",
1343 => x"00",
1344 => x"00",
1345 => x"00",
1346 => x"00",
1347 => x"00",
1348 => x"DC",
1349 => x"66",
1350 => x"66",
1351 => x"66",
1352 => x"7C",
1353 => x"60",
1354 => x"60",
1355 => x"F0",
1356 => x"00",
1357 => x"00",
1358 => x"00",
1359 => x"00",
1360 => x"76",
1361 => x"CC",
1362 => x"CC",
1363 => x"CC",
1364 => x"7C",
1365 => x"0C",
1366 => x"0C",
1367 => x"1E",
1368 => x"00",
1369 => x"00",
1370 => x"00",
1371 => x"00",
1372 => x"DC",
1373 => x"66",
1374 => x"60",
1375 => x"60",
1376 => x"60",
1377 => x"F0",
1378 => x"00",
1379 => x"00",
1380 => x"00",
1381 => x"00",
1382 => x"00",
1383 => x"00",
1384 => x"7C",
1385 => x"C6",
1386 => x"70",
1387 => x"1C",
1388 => x"C6",
1389 => x"7C",
1390 => x"00",
1391 => x"00",
1392 => x"00",
1393 => x"30",
1394 => x"30",
1395 => x"30",
1396 => x"FC",
1397 => x"30",
1398 => x"30",
1399 => x"30",
1400 => x"36",
1401 => x"1C",
1402 => x"00",
1403 => x"00",
1404 => x"00",
1405 => x"00",
1406 => x"00",
1407 => x"00",
1408 => x"CC",
1409 => x"CC",
1410 => x"CC",
1411 => x"CC",
1412 => x"CC",
1413 => x"76",
1414 => x"00",
1415 => x"00",
1416 => x"00",
1417 => x"00",
1418 => x"00",
1419 => x"00",
1420 => x"C6",
1421 => x"C6",
1422 => x"C6",
1423 => x"6C",
1424 => x"38",
1425 => x"10",
1426 => x"00",
1427 => x"00",
1428 => x"00",
1429 => x"00",
1430 => x"00",
1431 => x"00",
1432 => x"C6",
1433 => x"C6",
1434 => x"D6",
1435 => x"D6",
1436 => x"FE",
1437 => x"6C",
1438 => x"00",
1439 => x"00",
1440 => x"00",
1441 => x"00",
1442 => x"00",
1443 => x"00",
1444 => x"C6",
1445 => x"6C",
1446 => x"38",
1447 => x"38",
1448 => x"6C",
1449 => x"C6",
1450 => x"00",
1451 => x"00",
1452 => x"00",
1453 => x"00",
1454 => x"00",
1455 => x"00",
1456 => x"C6",
1457 => x"C6",
1458 => x"C6",
1459 => x"CE",
1460 => x"76",
1461 => x"06",
1462 => x"C6",
1463 => x"7C",
1464 => x"00",
1465 => x"00",
1466 => x"00",
1467 => x"00",
1468 => x"FE",
1469 => x"8C",
1470 => x"18",
1471 => x"30",
1472 => x"62",
1473 => x"FE",
1474 => x"00",
1475 => x"00",
1476 => x"00",
1477 => x"0E",
1478 => x"18",
1479 => x"18",
1480 => x"18",
1481 => x"70",
1482 => x"18",
1483 => x"18",
1484 => x"18",
1485 => x"0E",
1486 => x"00",
1487 => x"00",
1488 => x"00",
1489 => x"18",
1490 => x"18",
1491 => x"18",
1492 => x"18",
1493 => x"18",
1494 => x"18",
1495 => x"18",
1496 => x"18",
1497 => x"18",
1498 => x"00",
1499 => x"00",
1500 => x"00",
1501 => x"70",
1502 => x"18",
1503 => x"18",
1504 => x"18",
1505 => x"0E",
1506 => x"18",
1507 => x"18",
1508 => x"18",
1509 => x"70",
1510 => x"00",
1511 => x"00",
1512 => x"00",
1513 => x"76",
1514 => x"DC",
1515 => x"00",
1516 => x"00",
1517 => x"00",
1518 => x"00",
1519 => x"00",
1520 => x"00",
1521 => x"00",
1522 => x"00",
1523 => x"00",
1524 => x"66",
1525 => x"66",
1526 => x"00",
1527 => x"66",
1528 => x"66",
1529 => x"66",
1530 => x"3C",
1531 => x"18",
1532 => x"18",
1533 => x"3C",
1534 => x"00",
1535 => x"00",
1536 => x"30",
1537 => x"18",
1538 => x"00",
1539 => x"38",
1540 => x"6C",
1541 => x"C6",
1542 => x"C6",
1543 => x"FE",
1544 => x"C6",
1545 => x"C6",
1546 => x"00",
1547 => x"00",
1548 => x"18",
1549 => x"30",
1550 => x"00",
1551 => x"38",
1552 => x"6C",
1553 => x"C6",
1554 => x"C6",
1555 => x"FE",
1556 => x"C6",
1557 => x"C6",
1558 => x"00",
1559 => x"00",
1560 => x"38",
1561 => x"6C",
1562 => x"38",
1563 => x"00",
1564 => x"7C",
1565 => x"C6",
1566 => x"C6",
1567 => x"FE",
1568 => x"C6",
1569 => x"C6",
1570 => x"00",
1571 => x"00",
1572 => x"76",
1573 => x"DC",
1574 => x"00",
1575 => x"38",
1576 => x"6C",
1577 => x"C6",
1578 => x"C6",
1579 => x"FE",
1580 => x"C6",
1581 => x"C6",
1582 => x"00",
1583 => x"00",
1584 => x"6C",
1585 => x"6C",
1586 => x"00",
1587 => x"38",
1588 => x"6C",
1589 => x"C6",
1590 => x"C6",
1591 => x"FE",
1592 => x"C6",
1593 => x"C6",
1594 => x"00",
1595 => x"00",
1596 => x"38",
1597 => x"6C",
1598 => x"38",
1599 => x"00",
1600 => x"7C",
1601 => x"C6",
1602 => x"C6",
1603 => x"FE",
1604 => x"C6",
1605 => x"C6",
1606 => x"00",
1607 => x"00",
1608 => x"7E",
1609 => x"D8",
1610 => x"D8",
1611 => x"D8",
1612 => x"D8",
1613 => x"FE",
1614 => x"D8",
1615 => x"D8",
1616 => x"D8",
1617 => x"DE",
1618 => x"00",
1619 => x"00",
1620 => x"00",
1621 => x"3C",
1622 => x"66",
1623 => x"C0",
1624 => x"C0",
1625 => x"C0",
1626 => x"C6",
1627 => x"66",
1628 => x"3C",
1629 => x"18",
1630 => x"CC",
1631 => x"38",
1632 => x"18",
1633 => x"0C",
1634 => x"00",
1635 => x"FE",
1636 => x"66",
1637 => x"60",
1638 => x"7C",
1639 => x"60",
1640 => x"66",
1641 => x"FE",
1642 => x"00",
1643 => x"00",
1644 => x"18",
1645 => x"30",
1646 => x"00",
1647 => x"FE",
1648 => x"66",
1649 => x"60",
1650 => x"7C",
1651 => x"60",
1652 => x"66",
1653 => x"FE",
1654 => x"00",
1655 => x"00",
1656 => x"38",
1657 => x"6C",
1658 => x"00",
1659 => x"FE",
1660 => x"66",
1661 => x"60",
1662 => x"7C",
1663 => x"60",
1664 => x"66",
1665 => x"FE",
1666 => x"00",
1667 => x"00",
1668 => x"6C",
1669 => x"6C",
1670 => x"00",
1671 => x"FE",
1672 => x"66",
1673 => x"60",
1674 => x"7C",
1675 => x"60",
1676 => x"66",
1677 => x"FE",
1678 => x"00",
1679 => x"00",
1680 => x"18",
1681 => x"0C",
1682 => x"00",
1683 => x"3C",
1684 => x"18",
1685 => x"18",
1686 => x"18",
1687 => x"18",
1688 => x"18",
1689 => x"3C",
1690 => x"00",
1691 => x"00",
1692 => x"18",
1693 => x"30",
1694 => x"00",
1695 => x"3C",
1696 => x"18",
1697 => x"18",
1698 => x"18",
1699 => x"18",
1700 => x"18",
1701 => x"3C",
1702 => x"00",
1703 => x"00",
1704 => x"3C",
1705 => x"66",
1706 => x"00",
1707 => x"3C",
1708 => x"18",
1709 => x"18",
1710 => x"18",
1711 => x"18",
1712 => x"18",
1713 => x"3C",
1714 => x"00",
1715 => x"00",
1716 => x"66",
1717 => x"66",
1718 => x"00",
1719 => x"3C",
1720 => x"18",
1721 => x"18",
1722 => x"18",
1723 => x"18",
1724 => x"18",
1725 => x"3C",
1726 => x"00",
1727 => x"00",
1728 => x"00",
1729 => x"F8",
1730 => x"6C",
1731 => x"66",
1732 => x"66",
1733 => x"F6",
1734 => x"66",
1735 => x"66",
1736 => x"6C",
1737 => x"F8",
1738 => x"00",
1739 => x"00",
1740 => x"76",
1741 => x"DC",
1742 => x"00",
1743 => x"C6",
1744 => x"E6",
1745 => x"F6",
1746 => x"DE",
1747 => x"CE",
1748 => x"C6",
1749 => x"C6",
1750 => x"00",
1751 => x"00",
1752 => x"30",
1753 => x"18",
1754 => x"00",
1755 => x"7C",
1756 => x"C6",
1757 => x"C6",
1758 => x"C6",
1759 => x"C6",
1760 => x"C6",
1761 => x"7C",
1762 => x"00",
1763 => x"00",
1764 => x"18",
1765 => x"30",
1766 => x"00",
1767 => x"7C",
1768 => x"C6",
1769 => x"C6",
1770 => x"C6",
1771 => x"C6",
1772 => x"C6",
1773 => x"7C",
1774 => x"00",
1775 => x"00",
1776 => x"38",
1777 => x"6C",
1778 => x"00",
1779 => x"7C",
1780 => x"C6",
1781 => x"C6",
1782 => x"C6",
1783 => x"C6",
1784 => x"C6",
1785 => x"7C",
1786 => x"00",
1787 => x"00",
1788 => x"76",
1789 => x"DC",
1790 => x"00",
1791 => x"7C",
1792 => x"C6",
1793 => x"C6",
1794 => x"C6",
1795 => x"C6",
1796 => x"C6",
1797 => x"7C",
1798 => x"00",
1799 => x"00",
1800 => x"6C",
1801 => x"6C",
1802 => x"00",
1803 => x"7C",
1804 => x"C6",
1805 => x"C6",
1806 => x"C6",
1807 => x"C6",
1808 => x"C6",
1809 => x"7C",
1810 => x"00",
1811 => x"00",
1812 => x"00",
1813 => x"00",
1814 => x"00",
1815 => x"00",
1816 => x"6C",
1817 => x"38",
1818 => x"38",
1819 => x"6C",
1820 => x"00",
1821 => x"00",
1822 => x"00",
1823 => x"00",
1824 => x"00",
1825 => x"7E",
1826 => x"C6",
1827 => x"CE",
1828 => x"DE",
1829 => x"D6",
1830 => x"F6",
1831 => x"E6",
1832 => x"C6",
1833 => x"FC",
1834 => x"00",
1835 => x"00",
1836 => x"30",
1837 => x"18",
1838 => x"00",
1839 => x"C6",
1840 => x"C6",
1841 => x"C6",
1842 => x"C6",
1843 => x"C6",
1844 => x"C6",
1845 => x"7C",
1846 => x"00",
1847 => x"00",
1848 => x"18",
1849 => x"30",
1850 => x"00",
1851 => x"C6",
1852 => x"C6",
1853 => x"C6",
1854 => x"C6",
1855 => x"C6",
1856 => x"C6",
1857 => x"7C",
1858 => x"00",
1859 => x"00",
1860 => x"38",
1861 => x"6C",
1862 => x"00",
1863 => x"C6",
1864 => x"C6",
1865 => x"C6",
1866 => x"C6",
1867 => x"C6",
1868 => x"C6",
1869 => x"7C",
1870 => x"00",
1871 => x"00",
1872 => x"6C",
1873 => x"6C",
1874 => x"00",
1875 => x"C6",
1876 => x"C6",
1877 => x"C6",
1878 => x"C6",
1879 => x"C6",
1880 => x"C6",
1881 => x"7C",
1882 => x"00",
1883 => x"00",
1884 => x"0C",
1885 => x"18",
1886 => x"00",
1887 => x"66",
1888 => x"66",
1889 => x"66",
1890 => x"3C",
1891 => x"18",
1892 => x"18",
1893 => x"3C",
1894 => x"00",
1895 => x"00",
1896 => x"00",
1897 => x"F0",
1898 => x"60",
1899 => x"7C",
1900 => x"66",
1901 => x"66",
1902 => x"66",
1903 => x"7C",
1904 => x"60",
1905 => x"F0",
1906 => x"00",
1907 => x"00",
1908 => x"00",
1909 => x"7C",
1910 => x"C6",
1911 => x"C6",
1912 => x"C6",
1913 => x"CC",
1914 => x"C6",
1915 => x"C6",
1916 => x"D6",
1917 => x"DC",
1918 => x"80",
1919 => x"00",
1920 => x"00",
1921 => x"00",
1922 => x"00",
1923 => x"00",
1924 => x"00",
1925 => x"00",
1926 => x"00",
1927 => x"00",
1928 => x"00",
1929 => x"82",
1930 => x"FE",
1931 => x"00",
1932 => x"00",
1933 => x"00",
1934 => x"00",
1935 => x"18",
1936 => x"18",
1937 => x"00",
1938 => x"18",
1939 => x"18",
1940 => x"3C",
1941 => x"3C",
1942 => x"3C",
1943 => x"18",
1944 => x"00",
1945 => x"00",
1946 => x"10",
1947 => x"7C",
1948 => x"D6",
1949 => x"D0",
1950 => x"D0",
1951 => x"D6",
1952 => x"7C",
1953 => x"10",
1954 => x"00",
1955 => x"00",
1956 => x"00",
1957 => x"38",
1958 => x"6C",
1959 => x"60",
1960 => x"60",
1961 => x"F0",
1962 => x"60",
1963 => x"66",
1964 => x"F6",
1965 => x"6C",
1966 => x"00",
1967 => x"00",
1968 => x"00",
1969 => x"3C",
1970 => x"62",
1971 => x"60",
1972 => x"F8",
1973 => x"60",
1974 => x"F8",
1975 => x"60",
1976 => x"62",
1977 => x"3C",
1978 => x"00",
1979 => x"00",
1980 => x"00",
1981 => x"66",
1982 => x"66",
1983 => x"3C",
1984 => x"18",
1985 => x"7E",
1986 => x"18",
1987 => x"3C",
1988 => x"18",
1989 => x"18",
1990 => x"00",
1991 => x"00",
1992 => x"6C",
1993 => x"38",
1994 => x"00",
1995 => x"7C",
1996 => x"C6",
1997 => x"C0",
1998 => x"7C",
1999 => x"06",
2000 => x"C6",
2001 => x"7C",
2002 => x"00",
2003 => x"00",
2004 => x"7C",
2005 => x"C6",
2006 => x"C6",
2007 => x"60",
2008 => x"7C",
2009 => x"C6",
2010 => x"C6",
2011 => x"7C",
2012 => x"0C",
2013 => x"C6",
2014 => x"C6",
2015 => x"7C",
2016 => x"00",
2017 => x"6C",
2018 => x"38",
2019 => x"00",
2020 => x"7C",
2021 => x"C6",
2022 => x"70",
2023 => x"1C",
2024 => x"C6",
2025 => x"7C",
2026 => x"00",
2027 => x"00",
2028 => x"7E",
2029 => x"81",
2030 => x"99",
2031 => x"A5",
2032 => x"A1",
2033 => x"A1",
2034 => x"A5",
2035 => x"99",
2036 => x"81",
2037 => x"7E",
2038 => x"00",
2039 => x"00",
2040 => x"3C",
2041 => x"6C",
2042 => x"6C",
2043 => x"3E",
2044 => x"00",
2045 => x"7E",
2046 => x"00",
2047 => x"00",
2048 => x"00",
2049 => x"00",
2050 => x"00",
2051 => x"00",
2052 => x"00",
2053 => x"00",
2054 => x"00",
2055 => x"36",
2056 => x"6C",
2057 => x"D8",
2058 => x"6C",
2059 => x"36",
2060 => x"00",
2061 => x"00",
2062 => x"00",
2063 => x"00",
2064 => x"00",
2065 => x"00",
2066 => x"00",
2067 => x"00",
2068 => x"00",
2069 => x"7E",
2070 => x"06",
2071 => x"06",
2072 => x"06",
2073 => x"00",
2074 => x"00",
2075 => x"00",
2076 => x"00",
2077 => x"00",
2078 => x"00",
2079 => x"00",
2080 => x"00",
2081 => x"7E",
2082 => x"00",
2083 => x"00",
2084 => x"00",
2085 => x"00",
2086 => x"00",
2087 => x"00",
2088 => x"7E",
2089 => x"81",
2090 => x"B9",
2091 => x"A5",
2092 => x"A5",
2093 => x"B9",
2094 => x"A5",
2095 => x"A5",
2096 => x"81",
2097 => x"7E",
2098 => x"00",
2099 => x"00",
2100 => x"FF",
2101 => x"00",
2102 => x"00",
2103 => x"00",
2104 => x"00",
2105 => x"00",
2106 => x"00",
2107 => x"00",
2108 => x"00",
2109 => x"00",
2110 => x"00",
2111 => x"00",
2112 => x"00",
2113 => x"38",
2114 => x"6C",
2115 => x"38",
2116 => x"00",
2117 => x"00",
2118 => x"00",
2119 => x"00",
2120 => x"00",
2121 => x"00",
2122 => x"00",
2123 => x"00",
2124 => x"00",
2125 => x"00",
2126 => x"00",
2127 => x"18",
2128 => x"18",
2129 => x"7E",
2130 => x"18",
2131 => x"18",
2132 => x"00",
2133 => x"7E",
2134 => x"00",
2135 => x"00",
2136 => x"00",
2137 => x"38",
2138 => x"6C",
2139 => x"18",
2140 => x"30",
2141 => x"7C",
2142 => x"00",
2143 => x"00",
2144 => x"00",
2145 => x"00",
2146 => x"00",
2147 => x"00",
2148 => x"00",
2149 => x"38",
2150 => x"6C",
2151 => x"18",
2152 => x"6C",
2153 => x"38",
2154 => x"00",
2155 => x"00",
2156 => x"00",
2157 => x"00",
2158 => x"00",
2159 => x"00",
2160 => x"6C",
2161 => x"38",
2162 => x"00",
2163 => x"FE",
2164 => x"C6",
2165 => x"0C",
2166 => x"38",
2167 => x"62",
2168 => x"C6",
2169 => x"FE",
2170 => x"00",
2171 => x"00",
2172 => x"00",
2173 => x"00",
2174 => x"00",
2175 => x"00",
2176 => x"CC",
2177 => x"CC",
2178 => x"CC",
2179 => x"CC",
2180 => x"CC",
2181 => x"F6",
2182 => x"C0",
2183 => x"C0",
2184 => x"00",
2185 => x"7F",
2186 => x"DB",
2187 => x"DB",
2188 => x"DB",
2189 => x"7B",
2190 => x"1B",
2191 => x"1B",
2192 => x"1B",
2193 => x"1B",
2194 => x"00",
2195 => x"00",
2196 => x"00",
2197 => x"00",
2198 => x"00",
2199 => x"00",
2200 => x"00",
2201 => x"18",
2202 => x"18",
2203 => x"00",
2204 => x"00",
2205 => x"00",
2206 => x"00",
2207 => x"00",
2208 => x"00",
2209 => x"6C",
2210 => x"38",
2211 => x"00",
2212 => x"FE",
2213 => x"8C",
2214 => x"18",
2215 => x"30",
2216 => x"62",
2217 => x"FE",
2218 => x"00",
2219 => x"00",
2220 => x"00",
2221 => x"30",
2222 => x"70",
2223 => x"30",
2224 => x"30",
2225 => x"78",
2226 => x"00",
2227 => x"00",
2228 => x"00",
2229 => x"00",
2230 => x"00",
2231 => x"00",
2232 => x"38",
2233 => x"6C",
2234 => x"6C",
2235 => x"38",
2236 => x"00",
2237 => x"7C",
2238 => x"00",
2239 => x"00",
2240 => x"00",
2241 => x"00",
2242 => x"00",
2243 => x"00",
2244 => x"00",
2245 => x"00",
2246 => x"00",
2247 => x"D8",
2248 => x"6C",
2249 => x"36",
2250 => x"6C",
2251 => x"D8",
2252 => x"00",
2253 => x"00",
2254 => x"00",
2255 => x"00",
2256 => x"00",
2257 => x"6E",
2258 => x"DB",
2259 => x"DB",
2260 => x"DF",
2261 => x"D8",
2262 => x"D8",
2263 => x"D9",
2264 => x"DF",
2265 => x"6E",
2266 => x"00",
2267 => x"00",
2268 => x"00",
2269 => x"00",
2270 => x"00",
2271 => x"00",
2272 => x"6C",
2273 => x"DA",
2274 => x"DE",
2275 => x"D8",
2276 => x"DA",
2277 => x"6C",
2278 => x"00",
2279 => x"00",
2280 => x"66",
2281 => x"66",
2282 => x"00",
2283 => x"66",
2284 => x"66",
2285 => x"3C",
2286 => x"18",
2287 => x"18",
2288 => x"18",
2289 => x"3C",
2290 => x"00",
2291 => x"00",
2292 => x"00",
2293 => x"00",
2294 => x"00",
2295 => x"30",
2296 => x"30",
2297 => x"00",
2298 => x"30",
2299 => x"30",
2300 => x"60",
2301 => x"C6",
2302 => x"C6",
2303 => x"7C",
2304 => x"00",
2305 => x"00",
2306 => x"FF",
2307 => x"00",
2308 => x"00",
2309 => x"00",
2310 => x"00",
2311 => x"00",
2312 => x"00",
2313 => x"00",
2314 => x"00",
2315 => x"00",
2316 => x"18",
2317 => x"18",
2318 => x"18",
2319 => x"18",
2320 => x"18",
2321 => x"18",
2322 => x"00",
2323 => x"00",
2324 => x"00",
2325 => x"00",
2326 => x"00",
2327 => x"00",
2328 => x"00",
2329 => x"00",
2330 => x"00",
2331 => x"00",
2332 => x"00",
2333 => x"1F",
2334 => x"00",
2335 => x"00",
2336 => x"00",
2337 => x"00",
2338 => x"00",
2339 => x"00",
2340 => x"18",
2341 => x"18",
2342 => x"18",
2343 => x"18",
2344 => x"18",
2345 => x"1F",
2346 => x"00",
2347 => x"00",
2348 => x"00",
2349 => x"00",
2350 => x"00",
2351 => x"00",
2352 => x"00",
2353 => x"00",
2354 => x"00",
2355 => x"00",
2356 => x"00",
2357 => x"18",
2358 => x"18",
2359 => x"18",
2360 => x"18",
2361 => x"18",
2362 => x"18",
2363 => x"18",
2364 => x"18",
2365 => x"18",
2366 => x"18",
2367 => x"18",
2368 => x"18",
2369 => x"18",
2370 => x"18",
2371 => x"18",
2372 => x"18",
2373 => x"18",
2374 => x"18",
2375 => x"18",
2376 => x"00",
2377 => x"00",
2378 => x"00",
2379 => x"00",
2380 => x"00",
2381 => x"1F",
2382 => x"18",
2383 => x"18",
2384 => x"18",
2385 => x"18",
2386 => x"18",
2387 => x"18",
2388 => x"18",
2389 => x"18",
2390 => x"18",
2391 => x"18",
2392 => x"18",
2393 => x"1F",
2394 => x"18",
2395 => x"18",
2396 => x"18",
2397 => x"18",
2398 => x"18",
2399 => x"18",
2400 => x"00",
2401 => x"00",
2402 => x"00",
2403 => x"00",
2404 => x"00",
2405 => x"F8",
2406 => x"00",
2407 => x"00",
2408 => x"00",
2409 => x"00",
2410 => x"00",
2411 => x"00",
2412 => x"18",
2413 => x"18",
2414 => x"18",
2415 => x"18",
2416 => x"18",
2417 => x"F8",
2418 => x"00",
2419 => x"00",
2420 => x"00",
2421 => x"00",
2422 => x"00",
2423 => x"00",
2424 => x"00",
2425 => x"00",
2426 => x"00",
2427 => x"00",
2428 => x"00",
2429 => x"FF",
2430 => x"00",
2431 => x"00",
2432 => x"00",
2433 => x"00",
2434 => x"00",
2435 => x"00",
2436 => x"18",
2437 => x"18",
2438 => x"18",
2439 => x"18",
2440 => x"18",
2441 => x"FF",
2442 => x"00",
2443 => x"00",
2444 => x"00",
2445 => x"00",
2446 => x"00",
2447 => x"00",
2448 => x"00",
2449 => x"00",
2450 => x"00",
2451 => x"00",
2452 => x"00",
2453 => x"F8",
2454 => x"18",
2455 => x"18",
2456 => x"18",
2457 => x"18",
2458 => x"18",
2459 => x"18",
2460 => x"18",
2461 => x"18",
2462 => x"18",
2463 => x"18",
2464 => x"18",
2465 => x"F8",
2466 => x"18",
2467 => x"18",
2468 => x"18",
2469 => x"18",
2470 => x"18",
2471 => x"18",
2472 => x"00",
2473 => x"00",
2474 => x"00",
2475 => x"00",
2476 => x"00",
2477 => x"FF",
2478 => x"18",
2479 => x"18",
2480 => x"18",
2481 => x"18",
2482 => x"18",
2483 => x"18",
2484 => x"18",
2485 => x"18",
2486 => x"18",
2487 => x"18",
2488 => x"18",
2489 => x"FF",
2490 => x"18",
2491 => x"18",
2492 => x"18",
2493 => x"18",
2494 => x"18",
2495 => x"18",
2496 => x"00",
2497 => x"00",
2498 => x"00",
2499 => x"00",
2500 => x"00",
2501 => x"00",
2502 => x"00",
2503 => x"FF",
2504 => x"00",
2505 => x"00",
2506 => x"00",
2507 => x"00",
2508 => x"6C",
2509 => x"6C",
2510 => x"6C",
2511 => x"6C",
2512 => x"6C",
2513 => x"6C",
2514 => x"7C",
2515 => x"00",
2516 => x"00",
2517 => x"00",
2518 => x"00",
2519 => x"00",
2520 => x"00",
2521 => x"00",
2522 => x"00",
2523 => x"00",
2524 => x"3F",
2525 => x"30",
2526 => x"3F",
2527 => x"00",
2528 => x"00",
2529 => x"00",
2530 => x"00",
2531 => x"00",
2532 => x"6C",
2533 => x"6C",
2534 => x"6C",
2535 => x"6C",
2536 => x"6F",
2537 => x"60",
2538 => x"7F",
2539 => x"00",
2540 => x"00",
2541 => x"00",
2542 => x"00",
2543 => x"00",
2544 => x"00",
2545 => x"00",
2546 => x"00",
2547 => x"00",
2548 => x"7C",
2549 => x"6C",
2550 => x"6C",
2551 => x"6C",
2552 => x"6C",
2553 => x"6C",
2554 => x"6C",
2555 => x"6C",
2556 => x"6C",
2557 => x"6C",
2558 => x"6C",
2559 => x"6C",
2560 => x"6C",
2561 => x"6C",
2562 => x"6C",
2563 => x"6C",
2564 => x"6C",
2565 => x"6C",
2566 => x"6C",
2567 => x"6C",
2568 => x"00",
2569 => x"00",
2570 => x"00",
2571 => x"00",
2572 => x"7F",
2573 => x"60",
2574 => x"6F",
2575 => x"6C",
2576 => x"6C",
2577 => x"6C",
2578 => x"6C",
2579 => x"6C",
2580 => x"6C",
2581 => x"6C",
2582 => x"6C",
2583 => x"6C",
2584 => x"6F",
2585 => x"60",
2586 => x"6F",
2587 => x"6C",
2588 => x"6C",
2589 => x"6C",
2590 => x"6C",
2591 => x"6C",
2592 => x"00",
2593 => x"00",
2594 => x"00",
2595 => x"00",
2596 => x"FC",
2597 => x"0C",
2598 => x"FC",
2599 => x"00",
2600 => x"00",
2601 => x"00",
2602 => x"00",
2603 => x"00",
2604 => x"6C",
2605 => x"6C",
2606 => x"6C",
2607 => x"6C",
2608 => x"EC",
2609 => x"0C",
2610 => x"FC",
2611 => x"00",
2612 => x"00",
2613 => x"00",
2614 => x"00",
2615 => x"00",
2616 => x"00",
2617 => x"00",
2618 => x"00",
2619 => x"00",
2620 => x"FF",
2621 => x"00",
2622 => x"FF",
2623 => x"00",
2624 => x"00",
2625 => x"00",
2626 => x"00",
2627 => x"00",
2628 => x"6C",
2629 => x"6C",
2630 => x"6C",
2631 => x"6C",
2632 => x"EF",
2633 => x"00",
2634 => x"FF",
2635 => x"00",
2636 => x"00",
2637 => x"00",
2638 => x"00",
2639 => x"00",
2640 => x"00",
2641 => x"00",
2642 => x"00",
2643 => x"00",
2644 => x"FC",
2645 => x"0C",
2646 => x"EC",
2647 => x"6C",
2648 => x"6C",
2649 => x"6C",
2650 => x"6C",
2651 => x"6C",
2652 => x"6C",
2653 => x"6C",
2654 => x"6C",
2655 => x"6C",
2656 => x"EC",
2657 => x"0C",
2658 => x"EC",
2659 => x"6C",
2660 => x"6C",
2661 => x"6C",
2662 => x"6C",
2663 => x"6C",
2664 => x"00",
2665 => x"00",
2666 => x"00",
2667 => x"00",
2668 => x"FF",
2669 => x"00",
2670 => x"EF",
2671 => x"6C",
2672 => x"6C",
2673 => x"6C",
2674 => x"6C",
2675 => x"6C",
2676 => x"6C",
2677 => x"6C",
2678 => x"6C",
2679 => x"6C",
2680 => x"EF",
2681 => x"00",
2682 => x"EF",
2683 => x"6C",
2684 => x"6C",
2685 => x"6C",
2686 => x"6C",
2687 => x"6C",
2688 => x"60",
2689 => x"30",
2690 => x"18",
2691 => x"00",
2692 => x"78",
2693 => x"0C",
2694 => x"7C",
2695 => x"CC",
2696 => x"DC",
2697 => x"76",
2698 => x"00",
2699 => x"00",
2700 => x"18",
2701 => x"30",
2702 => x"60",
2703 => x"00",
2704 => x"78",
2705 => x"0C",
2706 => x"7C",
2707 => x"CC",
2708 => x"DC",
2709 => x"76",
2710 => x"00",
2711 => x"00",
2712 => x"30",
2713 => x"78",
2714 => x"CC",
2715 => x"00",
2716 => x"78",
2717 => x"0C",
2718 => x"7C",
2719 => x"CC",
2720 => x"DC",
2721 => x"76",
2722 => x"00",
2723 => x"00",
2724 => x"00",
2725 => x"76",
2726 => x"DC",
2727 => x"00",
2728 => x"78",
2729 => x"0C",
2730 => x"7C",
2731 => x"CC",
2732 => x"DC",
2733 => x"76",
2734 => x"00",
2735 => x"00",
2736 => x"00",
2737 => x"6C",
2738 => x"6C",
2739 => x"00",
2740 => x"78",
2741 => x"0C",
2742 => x"7C",
2743 => x"CC",
2744 => x"DC",
2745 => x"76",
2746 => x"00",
2747 => x"00",
2748 => x"38",
2749 => x"6C",
2750 => x"38",
2751 => x"00",
2752 => x"78",
2753 => x"0C",
2754 => x"7C",
2755 => x"CC",
2756 => x"DC",
2757 => x"76",
2758 => x"00",
2759 => x"00",
2760 => x"00",
2761 => x"00",
2762 => x"00",
2763 => x"7E",
2764 => x"DB",
2765 => x"1B",
2766 => x"7F",
2767 => x"D8",
2768 => x"DB",
2769 => x"7E",
2770 => x"00",
2771 => x"00",
2772 => x"00",
2773 => x"00",
2774 => x"00",
2775 => x"7C",
2776 => x"C6",
2777 => x"C0",
2778 => x"C0",
2779 => x"C6",
2780 => x"7C",
2781 => x"18",
2782 => x"6C",
2783 => x"38",
2784 => x"30",
2785 => x"18",
2786 => x"0C",
2787 => x"00",
2788 => x"7C",
2789 => x"C6",
2790 => x"FE",
2791 => x"C0",
2792 => x"C6",
2793 => x"7C",
2794 => x"00",
2795 => x"00",
2796 => x"0C",
2797 => x"18",
2798 => x"30",
2799 => x"00",
2800 => x"7C",
2801 => x"C6",
2802 => x"FE",
2803 => x"C0",
2804 => x"C6",
2805 => x"7C",
2806 => x"00",
2807 => x"00",
2808 => x"10",
2809 => x"38",
2810 => x"6C",
2811 => x"00",
2812 => x"7C",
2813 => x"C6",
2814 => x"FE",
2815 => x"C0",
2816 => x"C6",
2817 => x"7C",
2818 => x"00",
2819 => x"00",
2820 => x"00",
2821 => x"6C",
2822 => x"6C",
2823 => x"00",
2824 => x"7C",
2825 => x"C6",
2826 => x"FE",
2827 => x"C0",
2828 => x"C6",
2829 => x"7C",
2830 => x"00",
2831 => x"00",
2832 => x"60",
2833 => x"30",
2834 => x"18",
2835 => x"00",
2836 => x"38",
2837 => x"18",
2838 => x"18",
2839 => x"18",
2840 => x"18",
2841 => x"3C",
2842 => x"00",
2843 => x"00",
2844 => x"0C",
2845 => x"18",
2846 => x"30",
2847 => x"00",
2848 => x"38",
2849 => x"18",
2850 => x"18",
2851 => x"18",
2852 => x"18",
2853 => x"3C",
2854 => x"00",
2855 => x"00",
2856 => x"18",
2857 => x"3C",
2858 => x"66",
2859 => x"00",
2860 => x"38",
2861 => x"18",
2862 => x"18",
2863 => x"18",
2864 => x"18",
2865 => x"3C",
2866 => x"00",
2867 => x"00",
2868 => x"00",
2869 => x"6C",
2870 => x"6C",
2871 => x"00",
2872 => x"38",
2873 => x"18",
2874 => x"18",
2875 => x"18",
2876 => x"18",
2877 => x"3C",
2878 => x"00",
2879 => x"00",
2880 => x"78",
2881 => x"30",
2882 => x"78",
2883 => x"0C",
2884 => x"7E",
2885 => x"C6",
2886 => x"C6",
2887 => x"C6",
2888 => x"C6",
2889 => x"7C",
2890 => x"00",
2891 => x"00",
2892 => x"00",
2893 => x"76",
2894 => x"DC",
2895 => x"00",
2896 => x"DC",
2897 => x"66",
2898 => x"66",
2899 => x"66",
2900 => x"66",
2901 => x"66",
2902 => x"00",
2903 => x"00",
2904 => x"60",
2905 => x"30",
2906 => x"18",
2907 => x"00",
2908 => x"7C",
2909 => x"C6",
2910 => x"C6",
2911 => x"C6",
2912 => x"C6",
2913 => x"7C",
2914 => x"00",
2915 => x"00",
2916 => x"0C",
2917 => x"18",
2918 => x"30",
2919 => x"00",
2920 => x"7C",
2921 => x"C6",
2922 => x"C6",
2923 => x"C6",
2924 => x"C6",
2925 => x"7C",
2926 => x"00",
2927 => x"00",
2928 => x"10",
2929 => x"38",
2930 => x"6C",
2931 => x"00",
2932 => x"7C",
2933 => x"C6",
2934 => x"C6",
2935 => x"C6",
2936 => x"C6",
2937 => x"7C",
2938 => x"00",
2939 => x"00",
2940 => x"00",
2941 => x"76",
2942 => x"DC",
2943 => x"00",
2944 => x"7C",
2945 => x"C6",
2946 => x"C6",
2947 => x"C6",
2948 => x"C6",
2949 => x"7C",
2950 => x"00",
2951 => x"00",
2952 => x"00",
2953 => x"6C",
2954 => x"6C",
2955 => x"00",
2956 => x"7C",
2957 => x"C6",
2958 => x"C6",
2959 => x"C6",
2960 => x"C6",
2961 => x"7C",
2962 => x"00",
2963 => x"00",
2964 => x"00",
2965 => x"00",
2966 => x"18",
2967 => x"18",
2968 => x"00",
2969 => x"7E",
2970 => x"00",
2971 => x"18",
2972 => x"18",
2973 => x"00",
2974 => x"00",
2975 => x"00",
2976 => x"00",
2977 => x"00",
2978 => x"00",
2979 => x"00",
2980 => x"7E",
2981 => x"CE",
2982 => x"DE",
2983 => x"F6",
2984 => x"E6",
2985 => x"FC",
2986 => x"00",
2987 => x"00",
2988 => x"C0",
2989 => x"60",
2990 => x"30",
2991 => x"00",
2992 => x"CC",
2993 => x"CC",
2994 => x"CC",
2995 => x"CC",
2996 => x"CC",
2997 => x"76",
2998 => x"00",
2999 => x"00",
3000 => x"0C",
3001 => x"18",
3002 => x"30",
3003 => x"00",
3004 => x"CC",
3005 => x"CC",
3006 => x"CC",
3007 => x"CC",
3008 => x"CC",
3009 => x"76",
3010 => x"00",
3011 => x"00",
3012 => x"30",
3013 => x"78",
3014 => x"CC",
3015 => x"00",
3016 => x"CC",
3017 => x"CC",
3018 => x"CC",
3019 => x"CC",
3020 => x"CC",
3021 => x"76",
3022 => x"00",
3023 => x"00",
3024 => x"00",
3025 => x"CC",
3026 => x"CC",
3027 => x"00",
3028 => x"CC",
3029 => x"CC",
3030 => x"CC",
3031 => x"CC",
3032 => x"CC",
3033 => x"76",
3034 => x"00",
3035 => x"00",
3036 => x"0C",
3037 => x"18",
3038 => x"30",
3039 => x"00",
3040 => x"C6",
3041 => x"C6",
3042 => x"C6",
3043 => x"CE",
3044 => x"76",
3045 => x"06",
3046 => x"C6",
3047 => x"7C",
3048 => x"00",
3049 => x"F0",
3050 => x"60",
3051 => x"60",
3052 => x"78",
3053 => x"6C",
3054 => x"6C",
3055 => x"6C",
3056 => x"78",
3057 => x"60",
3058 => x"60",
3059 => x"F0",
3060 => x"00",
3061 => x"C6",
3062 => x"C6",
3063 => x"00",
3064 => x"C6",
3065 => x"C6",
3066 => x"C6",
3067 => x"CE",
3068 => x"76",
3069 => x"06",
3070 => x"C6",
3071 => x"7C",
others => X"42");
	attribute syn_ramstyle: string;
	attribute syn_ramstyle of mem: signal is "no_rw_check";
begin
	process (clka_i) -- Using port a.
	begin
	if (rising_edge(clka_i)) then
		if (wea_i = '1') then
		mem(conv_integer(addra_i)) <= dina_i;
			-- Using address bus a.
		end if;
		douta_o <= mem(conv_integer(addra_i));
	end if;
	end process;
	process (clkb_i) -- Using port b.
	begin
	if (rising_edge(clkb_i)) then
		if (web_i = '1') then
		mem(conv_integer(addrb_i)) <= dinb_i;
			-- Using address bus b.
		end if;
		doutb_o <= mem(conv_integer(addrb_i));
	end if;
	end process;
end rtl;
