-- from http://help.latticesemi.com/docs/webhelp/eng/wwhelp/wwhimpl/common/html/wwhelp.htm#href=Design%20Entry/inferring_ram_dual_port.htm
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
 
entity font_ub_dp_ram is
generic (
	addr_width : natural;
	data_width : natural);
port (
	addra_i	: in std_logic_vector (addr_width - 1 downto 0);
	wea_i	: in std_logic;
	clka_i	: in std_logic;
	dina_i	: in std_logic_vector (data_width - 1 downto 0);
	douta_o	: out std_logic_vector (data_width - 1 downto 0);
	addrb_i	: in std_logic_vector (addr_width - 1 downto 0);
	web_i	: in std_logic;
	clkb_i	: in std_logic;
	dinb_i	: in std_logic_vector (data_width - 1 downto 0);
	doutb_o	: out std_logic_vector (data_width - 1 downto 0));
end font_ub_dp_ram;
 
architecture rtl of font_ub_dp_ram is
	type mem_type is array ((2** addr_width) - 1 downto 0) of 
	std_logic_vector(data_width - 1 downto 0);
	signal mem : mem_type := (
-- even lines (upper byte)
-- char 0x00='\0' 
   0 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
   1 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
   2 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
   3 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x01='\x01
   4 =>	"01111110",	-- .######.
--   =>	"10000001",	-- #......#
   5 =>	"10100101",	-- #.#..#.#
--   =>	"10000001",	-- #......#
   6 =>	"10111101",	-- #.####.#
--   =>	"10011001",	-- #..##..#
   7 =>	"10000001",	-- #......#
--   =>	"01111110",	-- .######.

-- char 0x02='\x02
   8 =>	"01111110",	-- .######.
--   =>	"11111111",	-- ########
   9 =>	"11011011",	-- ##.##.##
--   =>	"11111111",	-- ########
  10 =>	"11000011",	-- ##....##
--   =>	"11100111",	-- ###..###
  11 =>	"11111111",	-- ########
--   =>	"01111110",	-- .######.

-- char 0x03='\x03
  12 =>	"01101100",	-- .##.##..
--   =>	"11111110",	-- #######.
  13 =>	"11111110",	-- #######.
--   =>	"11111110",	-- #######.
  14 =>	"01111100",	-- .#####..
--   =>	"00111000",	-- ..###...
  15 =>	"00010000",	-- ...#....
--   =>	"00000000",	-- ........

-- char 0x04='\x04
  16 =>	"00010000",	-- ...#....
--   =>	"00111000",	-- ..###...
  17 =>	"01111100",	-- .#####..
--   =>	"11111110",	-- #######.
  18 =>	"01111100",	-- .#####..
--   =>	"00111000",	-- ..###...
  19 =>	"00010000",	-- ...#....
--   =>	"00000000",	-- ........

-- char 0x05='\x05
  20 =>	"00111000",	-- ..###...
--   =>	"01111100",	-- .#####..
  21 =>	"00111000",	-- ..###...
--   =>	"11111110",	-- #######.
  22 =>	"11111110",	-- #######.
--   =>	"11010110",	-- ##.#.##.
  23 =>	"00010000",	-- ...#....
--   =>	"00111000",	-- ..###...

-- char 0x06='\x06
  24 =>	"00010000",	-- ...#....
--   =>	"00010000",	-- ...#....
  25 =>	"00111000",	-- ..###...
--   =>	"01111100",	-- .#####..
  26 =>	"11111110",	-- #######.
--   =>	"01111100",	-- .#####..
  27 =>	"00010000",	-- ...#....
--   =>	"00111000",	-- ..###...

-- char 0x07='\a' 
  28 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
  29 =>	"00011000",	-- ...##...
--   =>	"00111100",	-- ..####..
  30 =>	"00111100",	-- ..####..
--   =>	"00011000",	-- ...##...
  31 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x08='\b' 
  32 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
  33 =>	"11100111",	-- ###..###
--   =>	"11000011",	-- ##....##
  34 =>	"11000011",	-- ##....##
--   =>	"11100111",	-- ###..###
  35 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########

-- char 0x09='\t' 
  36 =>	"00000000",	-- ........
--   =>	"00111100",	-- ..####..
  37 =>	"01100110",	-- .##..##.
--   =>	"01000010",	-- .#....#.
  38 =>	"01000010",	-- .#....#.
--   =>	"01100110",	-- .##..##.
  39 =>	"00111100",	-- ..####..
--   =>	"00000000",	-- ........

-- char 0x0a='\n' 
  40 =>	"11111111",	-- ########
--   =>	"11000011",	-- ##....##
  41 =>	"10011001",	-- #..##..#
--   =>	"10111101",	-- #.####.#
  42 =>	"10111101",	-- #.####.#
--   =>	"10011001",	-- #..##..#
  43 =>	"11000011",	-- ##....##
--   =>	"11111111",	-- ########

-- char 0x0b='\v' 
  44 =>	"00001111",	-- ....####
--   =>	"00000111",	-- .....###
  45 =>	"00001111",	-- ....####
--   =>	"01111101",	-- .#####.#
  46 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
  47 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...

-- char 0x0c='\f' 
  48 =>	"00111100",	-- ..####..
--   =>	"01100110",	-- .##..##.
  49 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
  50 =>	"00111100",	-- ..####..
--   =>	"00011000",	-- ...##...
  51 =>	"01111110",	-- .######.
--   =>	"00011000",	-- ...##...

-- char 0x0d='\r' 
  52 =>	"00111111",	-- ..######
--   =>	"00110011",	-- ..##..##
  53 =>	"00111111",	-- ..######
--   =>	"00110000",	-- ..##....
  54 =>	"00110000",	-- ..##....
--   =>	"01110000",	-- .###....
  55 =>	"11110000",	-- ####....
--   =>	"11100000",	-- ###.....

-- char 0x0e='\x0e
  56 =>	"01111111",	-- .#######
--   =>	"01100011",	-- .##...##
  57 =>	"01111111",	-- .#######
--   =>	"01100011",	-- .##...##
  58 =>	"01100011",	-- .##...##
--   =>	"01100111",	-- .##..###
  59 =>	"11100110",	-- ###..##.
--   =>	"11000000",	-- ##......

-- char 0x0f='\x0f
  60 =>	"00011000",	-- ...##...
--   =>	"11011011",	-- ##.##.##
  61 =>	"00111100",	-- ..####..
--   =>	"11100111",	-- ###..###
  62 =>	"11100111",	-- ###..###
--   =>	"00111100",	-- ..####..
  63 =>	"11011011",	-- ##.##.##
--   =>	"00011000",	-- ...##...

-- char 0x10='\x10
  64 =>	"10000000",	-- #.......
--   =>	"11100000",	-- ###.....
  65 =>	"11111000",	-- #####...
--   =>	"11111110",	-- #######.
  66 =>	"11111000",	-- #####...
--   =>	"11100000",	-- ###.....
  67 =>	"10000000",	-- #.......
--   =>	"00000000",	-- ........

-- char 0x11='\x11
  68 =>	"00000010",	-- ......#.
--   =>	"00001110",	-- ....###.
  69 =>	"00111110",	-- ..#####.
--   =>	"11111110",	-- #######.
  70 =>	"00111110",	-- ..#####.
--   =>	"00001110",	-- ....###.
  71 =>	"00000010",	-- ......#.
--   =>	"00000000",	-- ........

-- char 0x12='\x12
  72 =>	"00011000",	-- ...##...
--   =>	"00111100",	-- ..####..
  73 =>	"01111110",	-- .######.
--   =>	"00011000",	-- ...##...
  74 =>	"00011000",	-- ...##...
--   =>	"01111110",	-- .######.
  75 =>	"00111100",	-- ..####..
--   =>	"00011000",	-- ...##...

-- char 0x13='\x13
  76 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
  77 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
  78 =>	"01100110",	-- .##..##.
--   =>	"00000000",	-- ........
  79 =>	"01100110",	-- .##..##.
--   =>	"00000000",	-- ........

-- char 0x14='\x14
  80 =>	"01111111",	-- .#######
--   =>	"11011011",	-- ##.##.##
  81 =>	"11011011",	-- ##.##.##
--   =>	"01111011",	-- .####.##
  82 =>	"00011011",	-- ...##.##
--   =>	"00011011",	-- ...##.##
  83 =>	"00011011",	-- ...##.##
--   =>	"00000000",	-- ........

-- char 0x15='\x15
  84 =>	"00111110",	-- ..#####.
--   =>	"01100011",	-- .##...##
  85 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
  86 =>	"01101100",	-- .##.##..
--   =>	"00111000",	-- ..###...
  87 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...

-- char 0x16='\x16
  88 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
  89 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
  90 =>	"01111110",	-- .######.
--   =>	"01111110",	-- .######.
  91 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........

-- char 0x17='\x17
  92 =>	"00011000",	-- ...##...
--   =>	"00111100",	-- ..####..
  93 =>	"01111110",	-- .######.
--   =>	"00011000",	-- ...##...
  94 =>	"01111110",	-- .######.
--   =>	"00111100",	-- ..####..
  95 =>	"00011000",	-- ...##...
--   =>	"11111111",	-- ########

-- char 0x18='\x18
  96 =>	"00011000",	-- ...##...
--   =>	"00111100",	-- ..####..
  97 =>	"01111110",	-- .######.
--   =>	"00011000",	-- ...##...
  98 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
  99 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........

-- char 0x19='\x19
 100 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 101 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 102 =>	"01111110",	-- .######.
--   =>	"00111100",	-- ..####..
 103 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........

-- char 0x1a='\x1a
 104 =>	"00000000",	-- ........
--   =>	"00011000",	-- ...##...
 105 =>	"00001100",	-- ....##..
--   =>	"11111110",	-- #######.
 106 =>	"00001100",	-- ....##..
--   =>	"00011000",	-- ...##...
 107 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x1b='\x1b
 108 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 109 =>	"01100000",	-- .##.....
--   =>	"11111110",	-- #######.
 110 =>	"01100000",	-- .##.....
--   =>	"00110000",	-- ..##....
 111 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x1c='\x1c
 112 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 113 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 114 =>	"11000000",	-- ##......
--   =>	"11111110",	-- #######.
 115 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x1d='\x1d
 116 =>	"00000000",	-- ........
--   =>	"00100100",	-- ..#..#..
 117 =>	"01100110",	-- .##..##.
--   =>	"11111111",	-- ########
 118 =>	"01100110",	-- .##..##.
--   =>	"00100100",	-- ..#..#..
 119 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x1e='\x1e
 120 =>	"00000000",	-- ........
--   =>	"00011000",	-- ...##...
 121 =>	"00111100",	-- ..####..
--   =>	"01111110",	-- .######.
 122 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 123 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x1f='\x1f
 124 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########
 125 =>	"11111111",	-- ########
--   =>	"01111110",	-- .######.
 126 =>	"00111100",	-- ..####..
--   =>	"00011000",	-- ...##...
 127 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x20=' '  
 128 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 129 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 130 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 131 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x21='!'  
 132 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 133 =>	"01111000",	-- .####...
--   =>	"00110000",	-- ..##....
 134 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 135 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........

-- char 0x22='\'' 
 136 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 137 =>	"01101100",	-- .##.##..
--   =>	"00000000",	-- ........
 138 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 139 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x23='#'  
 140 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 141 =>	"11111110",	-- #######.
--   =>	"01101100",	-- .##.##..
 142 =>	"11111110",	-- #######.
--   =>	"01101100",	-- .##.##..
 143 =>	"01101100",	-- .##.##..
--   =>	"00000000",	-- ........

-- char 0x24='$'  
 144 =>	"00110000",	-- ..##....
--   =>	"01111100",	-- .#####..
 145 =>	"11000000",	-- ##......
--   =>	"01111000",	-- .####...
 146 =>	"00001100",	-- ....##..
--   =>	"11111000",	-- #####...
 147 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........

-- char 0x25='%'  
 148 =>	"00000000",	-- ........
--   =>	"11000110",	-- ##...##.
 149 =>	"11001100",	-- ##..##..
--   =>	"00011000",	-- ...##...
 150 =>	"00110000",	-- ..##....
--   =>	"01100110",	-- .##..##.
 151 =>	"11000110",	-- ##...##.
--   =>	"00000000",	-- ........

-- char 0x26='&'  
 152 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 153 =>	"00111000",	-- ..###...
--   =>	"01110110",	-- .###.##.
 154 =>	"11011100",	-- ##.###..
--   =>	"11001100",	-- ##..##..
 155 =>	"01110110",	-- .###.##.
--   =>	"00000000",	-- ........

-- char 0x27='\"' 
 156 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 157 =>	"11000000",	-- ##......
--   =>	"00000000",	-- ........
 158 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 159 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x28='('  
 160 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
 161 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 162 =>	"01100000",	-- .##.....
--   =>	"00110000",	-- ..##....
 163 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........

-- char 0x29=')'  
 164 =>	"01100000",	-- .##.....
--   =>	"00110000",	-- ..##....
 165 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 166 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
 167 =>	"01100000",	-- .##.....
--   =>	"00000000",	-- ........

-- char 0x2a='*'  
 168 =>	"00000000",	-- ........
--   =>	"01100110",	-- .##..##.
 169 =>	"00111100",	-- ..####..
--   =>	"11111111",	-- ########
 170 =>	"00111100",	-- ..####..
--   =>	"01100110",	-- .##..##.
 171 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x2b='+'  
 172 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 173 =>	"00110000",	-- ..##....
--   =>	"11111100",	-- ######..
 174 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 175 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x2c=','  
 176 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 177 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 178 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 179 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....

-- char 0x2d='-'  
 180 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 181 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 182 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 183 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x2e='.'  
 184 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 185 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 186 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 187 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........

-- char 0x2f='/'  
 188 =>	"00000110",	-- .....##.
--   =>	"00001100",	-- ....##..
 189 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
 190 =>	"01100000",	-- .##.....
--   =>	"11000000",	-- ##......
 191 =>	"10000000",	-- #.......
--   =>	"00000000",	-- ........

-- char 0x30='0'  
 192 =>	"01111100",	-- .#####..
--   =>	"11000110",	-- ##...##.
 193 =>	"11001110",	-- ##..###.
--   =>	"11011110",	-- ##.####.
 194 =>	"11110110",	-- ####.##.
--   =>	"11100110",	-- ###..##.
 195 =>	"01111100",	-- .#####..
--   =>	"00000000",	-- ........

-- char 0x31='1'  
 196 =>	"00110000",	-- ..##....
--   =>	"01110000",	-- .###....
 197 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 198 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 199 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0x32='2'  
 200 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 201 =>	"00001100",	-- ....##..
--   =>	"00111000",	-- ..###...
 202 =>	"01100000",	-- .##.....
--   =>	"11001100",	-- ##..##..
 203 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0x33='3'  
 204 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 205 =>	"00001100",	-- ....##..
--   =>	"00111000",	-- ..###...
 206 =>	"00001100",	-- ....##..
--   =>	"11001100",	-- ##..##..
 207 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x34='4'  
 208 =>	"00011100",	-- ...###..
--   =>	"00111100",	-- ..####..
 209 =>	"01101100",	-- .##.##..
--   =>	"11001100",	-- ##..##..
 210 =>	"11111110",	-- #######.
--   =>	"00001100",	-- ....##..
 211 =>	"00011110",	-- ...####.
--   =>	"00000000",	-- ........

-- char 0x35='5'  
 212 =>	"11111100",	-- ######..
--   =>	"11000000",	-- ##......
 213 =>	"11111000",	-- #####...
--   =>	"00001100",	-- ....##..
 214 =>	"00001100",	-- ....##..
--   =>	"11001100",	-- ##..##..
 215 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x36='6'  
 216 =>	"00111000",	-- ..###...
--   =>	"01100000",	-- .##.....
 217 =>	"11000000",	-- ##......
--   =>	"11111000",	-- #####...
 218 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 219 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x37='7'  
 220 =>	"11111100",	-- ######..
--   =>	"11001100",	-- ##..##..
 221 =>	"00001100",	-- ....##..
--   =>	"00011000",	-- ...##...
 222 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 223 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........

-- char 0x38='8'  
 224 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 225 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 226 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 227 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x39='9'  
 228 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 229 =>	"11001100",	-- ##..##..
--   =>	"01111100",	-- .#####..
 230 =>	"00001100",	-- ....##..
--   =>	"00011000",	-- ...##...
 231 =>	"01110000",	-- .###....
--   =>	"00000000",	-- ........

-- char 0x3a=':'  
 232 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 233 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 234 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 235 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........

-- char 0x3b=';'  
 236 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 237 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 238 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 239 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....

-- char 0x3c='<'  
 240 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
 241 =>	"01100000",	-- .##.....
--   =>	"11000000",	-- ##......
 242 =>	"01100000",	-- .##.....
--   =>	"00110000",	-- ..##....
 243 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........

-- char 0x3d='='  
 244 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 245 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........
 246 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 247 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x3e='>'  
 248 =>	"01100000",	-- .##.....
--   =>	"00110000",	-- ..##....
 249 =>	"00011000",	-- ...##...
--   =>	"00001100",	-- ....##..
 250 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
 251 =>	"01100000",	-- .##.....
--   =>	"00000000",	-- ........

-- char 0x3f='?'  
 252 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 253 =>	"00001100",	-- ....##..
--   =>	"00011000",	-- ...##...
 254 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 255 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........

-- char 0x40='@'  
 256 =>	"01111100",	-- .#####..
--   =>	"11000110",	-- ##...##.
 257 =>	"11011110",	-- ##.####.
--   =>	"11011110",	-- ##.####.
 258 =>	"11011110",	-- ##.####.
--   =>	"11000000",	-- ##......
 259 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x41='A'  
 260 =>	"00110000",	-- ..##....
--   =>	"01111000",	-- .####...
 261 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 262 =>	"11111100",	-- ######..
--   =>	"11001100",	-- ##..##..
 263 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........

-- char 0x42='B'  
 264 =>	"11111100",	-- ######..
--   =>	"01100110",	-- .##..##.
 265 =>	"01100110",	-- .##..##.
--   =>	"01111100",	-- .#####..
 266 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 267 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0x43='C'  
 268 =>	"00111100",	-- ..####..
--   =>	"01100110",	-- .##..##.
 269 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 270 =>	"11000000",	-- ##......
--   =>	"01100110",	-- .##..##.
 271 =>	"00111100",	-- ..####..
--   =>	"00000000",	-- ........

-- char 0x44='D'  
 272 =>	"11111000",	-- #####...
--   =>	"01101100",	-- .##.##..
 273 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 274 =>	"01100110",	-- .##..##.
--   =>	"01101100",	-- .##.##..
 275 =>	"11111000",	-- #####...
--   =>	"00000000",	-- ........

-- char 0x45='E'  
 276 =>	"11111110",	-- #######.
--   =>	"01100010",	-- .##...#.
 277 =>	"01101000",	-- .##.#...
--   =>	"01111000",	-- .####...
 278 =>	"01101000",	-- .##.#...
--   =>	"01100010",	-- .##...#.
 279 =>	"11111110",	-- #######.
--   =>	"00000000",	-- ........

-- char 0x46='F'  
 280 =>	"11111110",	-- #######.
--   =>	"01100010",	-- .##...#.
 281 =>	"01101000",	-- .##.#...
--   =>	"01111000",	-- .####...
 282 =>	"01101000",	-- .##.#...
--   =>	"01100000",	-- .##.....
 283 =>	"11110000",	-- ####....
--   =>	"00000000",	-- ........

-- char 0x47='G'  
 284 =>	"00111100",	-- ..####..
--   =>	"01100110",	-- .##..##.
 285 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 286 =>	"11001110",	-- ##..###.
--   =>	"01100110",	-- .##..##.
 287 =>	"00111110",	-- ..#####.
--   =>	"00000000",	-- ........

-- char 0x48='H'  
 288 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 289 =>	"11001100",	-- ##..##..
--   =>	"11111100",	-- ######..
 290 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 291 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........

-- char 0x49='I'  
 292 =>	"01111000",	-- .####...
--   =>	"00110000",	-- ..##....
 293 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 294 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 295 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x4a='J'  
 296 =>	"00011110",	-- ...####.
--   =>	"00001100",	-- ....##..
 297 =>	"00001100",	-- ....##..
--   =>	"00001100",	-- ....##..
 298 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 299 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x4b='K'  
 300 =>	"11100110",	-- ###..##.
--   =>	"01100110",	-- .##..##.
 301 =>	"01101100",	-- .##.##..
--   =>	"01111000",	-- .####...
 302 =>	"01101100",	-- .##.##..
--   =>	"01100110",	-- .##..##.
 303 =>	"11100110",	-- ###..##.
--   =>	"00000000",	-- ........

-- char 0x4c='L'  
 304 =>	"11110000",	-- ####....
--   =>	"01100000",	-- .##.....
 305 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 306 =>	"01100010",	-- .##...#.
--   =>	"01100110",	-- .##..##.
 307 =>	"11111110",	-- #######.
--   =>	"00000000",	-- ........

-- char 0x4d='M'  
 308 =>	"11000110",	-- ##...##.
--   =>	"11101110",	-- ###.###.
 309 =>	"11111110",	-- #######.
--   =>	"11111110",	-- #######.
 310 =>	"11010110",	-- ##.#.##.
--   =>	"11000110",	-- ##...##.
 311 =>	"11000110",	-- ##...##.
--   =>	"00000000",	-- ........

-- char 0x4e='N'  
 312 =>	"11000110",	-- ##...##.
--   =>	"11100110",	-- ###..##.
 313 =>	"11110110",	-- ####.##.
--   =>	"11011110",	-- ##.####.
 314 =>	"11001110",	-- ##..###.
--   =>	"11000110",	-- ##...##.
 315 =>	"11000110",	-- ##...##.
--   =>	"00000000",	-- ........

-- char 0x4f='O'  
 316 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 317 =>	"11000110",	-- ##...##.
--   =>	"11000110",	-- ##...##.
 318 =>	"11000110",	-- ##...##.
--   =>	"01101100",	-- .##.##..
 319 =>	"00111000",	-- ..###...
--   =>	"00000000",	-- ........

-- char 0x50='P'  
 320 =>	"11111100",	-- ######..
--   =>	"01100110",	-- .##..##.
 321 =>	"01100110",	-- .##..##.
--   =>	"01111100",	-- .#####..
 322 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 323 =>	"11110000",	-- ####....
--   =>	"00000000",	-- ........

-- char 0x51='Q'  
 324 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 325 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 326 =>	"11011100",	-- ##.###..
--   =>	"01111000",	-- .####...
 327 =>	"00011100",	-- ...###..
--   =>	"00000000",	-- ........

-- char 0x52='R'  
 328 =>	"11111100",	-- ######..
--   =>	"01100110",	-- .##..##.
 329 =>	"01100110",	-- .##..##.
--   =>	"01111100",	-- .#####..
 330 =>	"01101100",	-- .##.##..
--   =>	"01100110",	-- .##..##.
 331 =>	"11100110",	-- ###..##.
--   =>	"00000000",	-- ........

-- char 0x53='S'  
 332 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 333 =>	"01100000",	-- .##.....
--   =>	"00110000",	-- ..##....
 334 =>	"00011000",	-- ...##...
--   =>	"11001100",	-- ##..##..
 335 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x54='T'  
 336 =>	"11111100",	-- ######..
--   =>	"10110100",	-- #.##.#..
 337 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 338 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 339 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x55='U'  
 340 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 341 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 342 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 343 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0x56='V'  
 344 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 345 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 346 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 347 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........

-- char 0x57='W'  
 348 =>	"11000110",	-- ##...##.
--   =>	"11000110",	-- ##...##.
 349 =>	"11000110",	-- ##...##.
--   =>	"11010110",	-- ##.#.##.
 350 =>	"11111110",	-- #######.
--   =>	"11101110",	-- ###.###.
 351 =>	"11000110",	-- ##...##.
--   =>	"00000000",	-- ........

-- char 0x58='X'  
 352 =>	"11000110",	-- ##...##.
--   =>	"11000110",	-- ##...##.
 353 =>	"01101100",	-- .##.##..
--   =>	"00111000",	-- ..###...
 354 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 355 =>	"11000110",	-- ##...##.
--   =>	"00000000",	-- ........

-- char 0x59='Y'  
 356 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 357 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 358 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 359 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x5a='Z'  
 360 =>	"11111110",	-- #######.
--   =>	"11000110",	-- ##...##.
 361 =>	"10001100",	-- #...##..
--   =>	"00011000",	-- ...##...
 362 =>	"00110010",	-- ..##..#.
--   =>	"01100110",	-- .##..##.
 363 =>	"11111110",	-- #######.
--   =>	"00000000",	-- ........

-- char 0x5b='['  
 364 =>	"01111000",	-- .####...
--   =>	"01100000",	-- .##.....
 365 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 366 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 367 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x5c='\\' 
 368 =>	"11000000",	-- ##......
--   =>	"01100000",	-- .##.....
 369 =>	"00110000",	-- ..##....
--   =>	"00011000",	-- ...##...
 370 =>	"00001100",	-- ....##..
--   =>	"00000110",	-- .....##.
 371 =>	"00000010",	-- ......#.
--   =>	"00000000",	-- ........

-- char 0x5d=']'  
 372 =>	"01111000",	-- .####...
--   =>	"00011000",	-- ...##...
 373 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 374 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 375 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x5e='^'  
 376 =>	"00010000",	-- ...#....
--   =>	"00111000",	-- ..###...
 377 =>	"01101100",	-- .##.##..
--   =>	"11000110",	-- ##...##.
 378 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 379 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x5f='_'  
 380 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 381 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 382 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 383 =>	"00000000",	-- ........
--   =>	"11111111",	-- ########

-- char 0x60='`'  
 384 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 385 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........
 386 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 387 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x61='a'  
 388 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 389 =>	"01111000",	-- .####...
--   =>	"00001100",	-- ....##..
 390 =>	"01111100",	-- .#####..
--   =>	"11001100",	-- ##..##..
 391 =>	"01110110",	-- .###.##.
--   =>	"00000000",	-- ........

-- char 0x62='b'  
 392 =>	"11100000",	-- ###.....
--   =>	"01100000",	-- .##.....
 393 =>	"01100000",	-- .##.....
--   =>	"01111100",	-- .#####..
 394 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 395 =>	"11011100",	-- ##.###..
--   =>	"00000000",	-- ........

-- char 0x63='c'  
 396 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 397 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 398 =>	"11000000",	-- ##......
--   =>	"11001100",	-- ##..##..
 399 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x64='d'  
 400 =>	"00011100",	-- ...###..
--   =>	"00001100",	-- ....##..
 401 =>	"00001100",	-- ....##..
--   =>	"01111100",	-- .#####..
 402 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 403 =>	"01110110",	-- .###.##.
--   =>	"00000000",	-- ........

-- char 0x65='e'  
 404 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 405 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 406 =>	"11111100",	-- ######..
--   =>	"11000000",	-- ##......
 407 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x66='f'  
 408 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 409 =>	"01100000",	-- .##.....
--   =>	"11110000",	-- ####....
 410 =>	"01100000",	-- .##.....
--   =>	"01100000",	-- .##.....
 411 =>	"11110000",	-- ####....
--   =>	"00000000",	-- ........

-- char 0x67='g'  
 412 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 413 =>	"01110110",	-- .###.##.
--   =>	"11001100",	-- ##..##..
 414 =>	"11001100",	-- ##..##..
--   =>	"01111100",	-- .#####..
 415 =>	"00001100",	-- ....##..
--   =>	"11111000",	-- #####...

-- char 0x68='h'  
 416 =>	"11100000",	-- ###.....
--   =>	"01100000",	-- .##.....
 417 =>	"01101100",	-- .##.##..
--   =>	"01110110",	-- .###.##.
 418 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 419 =>	"11100110",	-- ###..##.
--   =>	"00000000",	-- ........

-- char 0x69='i'  
 420 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 421 =>	"01110000",	-- .###....
--   =>	"00110000",	-- ..##....
 422 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 423 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x6a='j'  
 424 =>	"00001100",	-- ....##..
--   =>	"00000000",	-- ........
 425 =>	"00001100",	-- ....##..
--   =>	"00001100",	-- ....##..
 426 =>	"00001100",	-- ....##..
--   =>	"11001100",	-- ##..##..
 427 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...

-- char 0x6b='k'  
 428 =>	"11100000",	-- ###.....
--   =>	"01100000",	-- .##.....
 429 =>	"01100110",	-- .##..##.
--   =>	"01101100",	-- .##.##..
 430 =>	"01111000",	-- .####...
--   =>	"01101100",	-- .##.##..
 431 =>	"11100110",	-- ###..##.
--   =>	"00000000",	-- ........

-- char 0x6c='l'  
 432 =>	"01110000",	-- .###....
--   =>	"00110000",	-- ..##....
 433 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 434 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 435 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x6d='m'  
 436 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 437 =>	"11001100",	-- ##..##..
--   =>	"11111110",	-- #######.
 438 =>	"11111110",	-- #######.
--   =>	"11010110",	-- ##.#.##.
 439 =>	"11000110",	-- ##...##.
--   =>	"00000000",	-- ........

-- char 0x6e='n'  
 440 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 441 =>	"11111000",	-- #####...
--   =>	"11001100",	-- ##..##..
 442 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 443 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........

-- char 0x6f='o'  
 444 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 445 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 446 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 447 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x70='p'  
 448 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 449 =>	"11011100",	-- ##.###..
--   =>	"01100110",	-- .##..##.
 450 =>	"01100110",	-- .##..##.
--   =>	"01111100",	-- .#####..
 451 =>	"01100000",	-- .##.....
--   =>	"11110000",	-- ####....

-- char 0x71='q'  
 452 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 453 =>	"01110110",	-- .###.##.
--   =>	"11001100",	-- ##..##..
 454 =>	"11001100",	-- ##..##..
--   =>	"01111100",	-- .#####..
 455 =>	"00001100",	-- ....##..
--   =>	"00011110",	-- ...####.

-- char 0x72='r'  
 456 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 457 =>	"11011100",	-- ##.###..
--   =>	"01110110",	-- .###.##.
 458 =>	"01100110",	-- .##..##.
--   =>	"01100000",	-- .##.....
 459 =>	"11110000",	-- ####....
--   =>	"00000000",	-- ........

-- char 0x73='s'  
 460 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 461 =>	"01111100",	-- .#####..
--   =>	"11000000",	-- ##......
 462 =>	"01111000",	-- .####...
--   =>	"00001100",	-- ....##..
 463 =>	"11111000",	-- #####...
--   =>	"00000000",	-- ........

-- char 0x74='t'  
 464 =>	"00010000",	-- ...#....
--   =>	"00110000",	-- ..##....
 465 =>	"01111100",	-- .#####..
--   =>	"00110000",	-- ..##....
 466 =>	"00110000",	-- ..##....
--   =>	"00110100",	-- ..##.#..
 467 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........

-- char 0x75='u'  
 468 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 469 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 470 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 471 =>	"01110110",	-- .###.##.
--   =>	"00000000",	-- ........

-- char 0x76='v'  
 472 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 473 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 474 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 475 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........

-- char 0x77='w'  
 476 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 477 =>	"11000110",	-- ##...##.
--   =>	"11010110",	-- ##.#.##.
 478 =>	"11111110",	-- #######.
--   =>	"11111110",	-- #######.
 479 =>	"01101100",	-- .##.##..
--   =>	"00000000",	-- ........

-- char 0x78='x'  
 480 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 481 =>	"11000110",	-- ##...##.
--   =>	"01101100",	-- .##.##..
 482 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 483 =>	"11000110",	-- ##...##.
--   =>	"00000000",	-- ........

-- char 0x79='y'  
 484 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 485 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 486 =>	"11001100",	-- ##..##..
--   =>	"01111100",	-- .#####..
 487 =>	"00001100",	-- ....##..
--   =>	"11111000",	-- #####...

-- char 0x7a='z'  
 488 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 489 =>	"11111100",	-- ######..
--   =>	"10011000",	-- #..##...
 490 =>	"00110000",	-- ..##....
--   =>	"01100100",	-- .##..#..
 491 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0x7b='{'  
 492 =>	"00011100",	-- ...###..
--   =>	"00110000",	-- ..##....
 493 =>	"00110000",	-- ..##....
--   =>	"11100000",	-- ###.....
 494 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 495 =>	"00011100",	-- ...###..
--   =>	"00000000",	-- ........

-- char 0x7c='|'  
 496 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 497 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........
 498 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 499 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........

-- char 0x7d='}'  
 500 =>	"11100000",	-- ###.....
--   =>	"00110000",	-- ..##....
 501 =>	"00110000",	-- ..##....
--   =>	"00011100",	-- ...###..
 502 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 503 =>	"11100000",	-- ###.....
--   =>	"00000000",	-- ........

-- char 0x7e='~'  
 504 =>	"01110110",	-- .###.##.
--   =>	"11011100",	-- ##.###..
 505 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 506 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 507 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0x7f='\x7f
 508 =>	"00000000",	-- ........
--   =>	"00010000",	-- ...#....
 509 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 510 =>	"11000110",	-- ##...##.
--   =>	"11000110",	-- ##...##.
 511 =>	"11111110",	-- #######.
--   =>	"00000000",	-- ........

-- char 0x80='\x80
 512 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 513 =>	"11000000",	-- ##......
--   =>	"11001100",	-- ##..##..
 514 =>	"01111000",	-- .####...
--   =>	"00011000",	-- ...##...
 515 =>	"00001100",	-- ....##..
--   =>	"01111000",	-- .####...

-- char 0x81='\x81
 516 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 517 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 518 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 519 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........

-- char 0x82='\x82
 520 =>	"00011100",	-- ...###..
--   =>	"00000000",	-- ........
 521 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 522 =>	"11111100",	-- ######..
--   =>	"11000000",	-- ##......
 523 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x83='\x83
 524 =>	"01111110",	-- .######.
--   =>	"11000011",	-- ##....##
 525 =>	"00111100",	-- ..####..
--   =>	"00000110",	-- .....##.
 526 =>	"00111110",	-- ..#####.
--   =>	"01100110",	-- .##..##.
 527 =>	"00111111",	-- ..######
--   =>	"00000000",	-- ........

-- char 0x84='\x84
 528 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........
 529 =>	"01111000",	-- .####...
--   =>	"00001100",	-- ....##..
 530 =>	"01111100",	-- .#####..
--   =>	"11001100",	-- ##..##..
 531 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........

-- char 0x85='\x85
 532 =>	"11100000",	-- ###.....
--   =>	"00000000",	-- ........
 533 =>	"01111000",	-- .####...
--   =>	"00001100",	-- ....##..
 534 =>	"01111100",	-- .#####..
--   =>	"11001100",	-- ##..##..
 535 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........

-- char 0x86='\x86
 536 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 537 =>	"01111000",	-- .####...
--   =>	"00001100",	-- ....##..
 538 =>	"01111100",	-- .#####..
--   =>	"11001100",	-- ##..##..
 539 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........

-- char 0x87='\x87
 540 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 541 =>	"01111000",	-- .####...
--   =>	"11000000",	-- ##......
 542 =>	"11000000",	-- ##......
--   =>	"01111000",	-- .####...
 543 =>	"00001100",	-- ....##..
--   =>	"00111000",	-- ..###...

-- char 0x88='\x88
 544 =>	"01111110",	-- .######.
--   =>	"11000011",	-- ##....##
 545 =>	"00111100",	-- ..####..
--   =>	"01100110",	-- .##..##.
 546 =>	"01111110",	-- .######.
--   =>	"01100000",	-- .##.....
 547 =>	"00111100",	-- ..####..
--   =>	"00000000",	-- ........

-- char 0x89='\x89
 548 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........
 549 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 550 =>	"11111100",	-- ######..
--   =>	"11000000",	-- ##......
 551 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x8a='\x8a
 552 =>	"11100000",	-- ###.....
--   =>	"00000000",	-- ........
 553 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 554 =>	"11111100",	-- ######..
--   =>	"11000000",	-- ##......
 555 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x8b='\x8b
 556 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........
 557 =>	"01110000",	-- .###....
--   =>	"00110000",	-- ..##....
 558 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 559 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x8c='\x8c
 560 =>	"01111100",	-- .#####..
--   =>	"11000110",	-- ##...##.
 561 =>	"00111000",	-- ..###...
--   =>	"00011000",	-- ...##...
 562 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 563 =>	"00111100",	-- ..####..
--   =>	"00000000",	-- ........

-- char 0x8d='\x8d
 564 =>	"11100000",	-- ###.....
--   =>	"00000000",	-- ........
 565 =>	"01110000",	-- .###....
--   =>	"00110000",	-- ..##....
 566 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 567 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x8e='\x8e
 568 =>	"11000110",	-- ##...##.
--   =>	"00111000",	-- ..###...
 569 =>	"01101100",	-- .##.##..
--   =>	"11000110",	-- ##...##.
 570 =>	"11111110",	-- #######.
--   =>	"11000110",	-- ##...##.
 571 =>	"11000110",	-- ##...##.
--   =>	"00000000",	-- ........

-- char 0x8f='\x8f
 572 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 573 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 574 =>	"11001100",	-- ##..##..
--   =>	"11111100",	-- ######..
 575 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........

-- char 0x90='\x90
 576 =>	"00011100",	-- ...###..
--   =>	"00000000",	-- ........
 577 =>	"11111100",	-- ######..
--   =>	"01100000",	-- .##.....
 578 =>	"01111000",	-- .####...
--   =>	"01100000",	-- .##.....
 579 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0x91='\x91
 580 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 581 =>	"01111111",	-- .#######
--   =>	"00001100",	-- ....##..
 582 =>	"01111111",	-- .#######
--   =>	"11001100",	-- ##..##..
 583 =>	"01111111",	-- .#######
--   =>	"00000000",	-- ........

-- char 0x92='\x92
 584 =>	"00111110",	-- ..#####.
--   =>	"01101100",	-- .##.##..
 585 =>	"11001100",	-- ##..##..
--   =>	"11111110",	-- #######.
 586 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 587 =>	"11001110",	-- ##..###.
--   =>	"00000000",	-- ........

-- char 0x93='\x93
 588 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 589 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 590 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 591 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x94='\x94
 592 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 593 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 594 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 595 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x95='\x95
 596 =>	"00000000",	-- ........
--   =>	"11100000",	-- ###.....
 597 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 598 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 599 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x96='\x96
 600 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 601 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 602 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 603 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........

-- char 0x97='\x97
 604 =>	"00000000",	-- ........
--   =>	"11100000",	-- ###.....
 605 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 606 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 607 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........

-- char 0x98='\x98
 608 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 609 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 610 =>	"11001100",	-- ##..##..
--   =>	"01111100",	-- .#####..
 611 =>	"00001100",	-- ....##..
--   =>	"11111000",	-- #####...

-- char 0x99='\x99
 612 =>	"11000011",	-- ##....##
--   =>	"00011000",	-- ...##...
 613 =>	"00111100",	-- ..####..
--   =>	"01100110",	-- .##..##.
 614 =>	"01100110",	-- .##..##.
--   =>	"00111100",	-- ..####..
 615 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........

-- char 0x9a='\x9a
 616 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........
 617 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 618 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 619 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0x9b='\x9b
 620 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 621 =>	"01111110",	-- .######.
--   =>	"11000000",	-- ##......
 622 =>	"11000000",	-- ##......
--   =>	"01111110",	-- .######.
 623 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0x9c='\x9c
 624 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 625 =>	"01100100",	-- .##..#..
--   =>	"11110000",	-- ####....
 626 =>	"01100000",	-- .##.....
--   =>	"11100110",	-- ###..##.
 627 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0x9d='\x9d
 628 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 629 =>	"01111000",	-- .####...
--   =>	"11111100",	-- ######..
 630 =>	"00110000",	-- ..##....
--   =>	"11111100",	-- ######..
 631 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....

-- char 0x9e='\x9e
 632 =>	"11111000",	-- #####...
--   =>	"11001100",	-- ##..##..
 633 =>	"11001100",	-- ##..##..
--   =>	"11111010",	-- #####.#.
 634 =>	"11000110",	-- ##...##.
--   =>	"11001111",	-- ##..####
 635 =>	"11000110",	-- ##...##.
--   =>	"11000111",	-- ##...###

-- char 0x9f='\x9f
 636 =>	"00001110",	-- ....###.
--   =>	"00011011",	-- ...##.##
 637 =>	"00011000",	-- ...##...
--   =>	"00111100",	-- ..####..
 638 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 639 =>	"11011000",	-- ##.##...
--   =>	"01110000",	-- .###....

-- char 0xa0='\xa0
 640 =>	"00011100",	-- ...###..
--   =>	"00000000",	-- ........
 641 =>	"01111000",	-- .####...
--   =>	"00001100",	-- ....##..
 642 =>	"01111100",	-- .#####..
--   =>	"11001100",	-- ##..##..
 643 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........

-- char 0xa1='\xa1
 644 =>	"00111000",	-- ..###...
--   =>	"00000000",	-- ........
 645 =>	"01110000",	-- .###....
--   =>	"00110000",	-- ..##....
 646 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 647 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0xa2='\xa2
 648 =>	"00000000",	-- ........
--   =>	"00011100",	-- ...###..
 649 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 650 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 651 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0xa3='\xa3
 652 =>	"00000000",	-- ........
--   =>	"00011100",	-- ...###..
 653 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 654 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 655 =>	"01111110",	-- .######.
--   =>	"00000000",	-- ........

-- char 0xa4='\xa4
 656 =>	"00000000",	-- ........
--   =>	"11111000",	-- #####...
 657 =>	"00000000",	-- ........
--   =>	"11111000",	-- #####...
 658 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 659 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........

-- char 0xa5='\xa5
 660 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........
 661 =>	"11001100",	-- ##..##..
--   =>	"11101100",	-- ###.##..
 662 =>	"11111100",	-- ######..
--   =>	"11011100",	-- ##.###..
 663 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........

-- char 0xa6='\xa6
 664 =>	"00111100",	-- ..####..
--   =>	"01101100",	-- .##.##..
 665 =>	"01101100",	-- .##.##..
--   =>	"00111110",	-- ..#####.
 666 =>	"00000000",	-- ........
--   =>	"01111110",	-- .######.
 667 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xa7='\xa7
 668 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 669 =>	"01101100",	-- .##.##..
--   =>	"00111000",	-- ..###...
 670 =>	"00000000",	-- ........
--   =>	"01111100",	-- .#####..
 671 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xa8='\xa8
 672 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 673 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
 674 =>	"11000000",	-- ##......
--   =>	"11001100",	-- ##..##..
 675 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0xa9='\xa9
 676 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 677 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 678 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 679 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xaa='\xaa
 680 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 681 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 682 =>	"00001100",	-- ....##..
--   =>	"00001100",	-- ....##..
 683 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xab='\xab
 684 =>	"11000011",	-- ##....##
--   =>	"11000110",	-- ##...##.
 685 =>	"11001100",	-- ##..##..
--   =>	"11011110",	-- ##.####.
 686 =>	"00110011",	-- ..##..##
--   =>	"01100110",	-- .##..##.
 687 =>	"11001100",	-- ##..##..
--   =>	"00001111",	-- ....####

-- char 0xac='\xac
 688 =>	"11000011",	-- ##....##
--   =>	"11000110",	-- ##...##.
 689 =>	"11001100",	-- ##..##..
--   =>	"11011011",	-- ##.##.##
 690 =>	"00110111",	-- ..##.###
--   =>	"01101111",	-- .##.####
 691 =>	"11001111",	-- ##..####
--   =>	"00000011",	-- ......##

-- char 0xad='\xad
 692 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 693 =>	"00000000",	-- ........
--   =>	"00011000",	-- ...##...
 694 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 695 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........

-- char 0xae='\xae
 696 =>	"00000000",	-- ........
--   =>	"00110011",	-- ..##..##
 697 =>	"01100110",	-- .##..##.
--   =>	"11001100",	-- ##..##..
 698 =>	"01100110",	-- .##..##.
--   =>	"00110011",	-- ..##..##
 699 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xaf='\xaf
 700 =>	"00000000",	-- ........
--   =>	"11001100",	-- ##..##..
 701 =>	"01100110",	-- .##..##.
--   =>	"00110011",	-- ..##..##
 702 =>	"01100110",	-- .##..##.
--   =>	"11001100",	-- ##..##..
 703 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xb0='\xb0
 704 =>	"00100010",	-- ..#...#.
--   =>	"10001000",	-- #...#...
 705 =>	"00100010",	-- ..#...#.
--   =>	"10001000",	-- #...#...
 706 =>	"00100010",	-- ..#...#.
--   =>	"10001000",	-- #...#...
 707 =>	"00100010",	-- ..#...#.
--   =>	"10001000",	-- #...#...

-- char 0xb1='\xb1
 708 =>	"01010101",	-- .#.#.#.#
--   =>	"10101010",	-- #.#.#.#.
 709 =>	"01010101",	-- .#.#.#.#
--   =>	"10101010",	-- #.#.#.#.
 710 =>	"01010101",	-- .#.#.#.#
--   =>	"10101010",	-- #.#.#.#.
 711 =>	"01010101",	-- .#.#.#.#
--   =>	"10101010",	-- #.#.#.#.

-- char 0xb2='\xb2
 712 =>	"11011011",	-- ##.##.##
--   =>	"01110111",	-- .###.###
 713 =>	"11011011",	-- ##.##.##
--   =>	"11101110",	-- ###.###.
 714 =>	"11011011",	-- ##.##.##
--   =>	"01110111",	-- .###.###
 715 =>	"11011011",	-- ##.##.##
--   =>	"11101110",	-- ###.###.

-- char 0xb3='\xb3
 716 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 717 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 718 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 719 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xb4='\xb4
 720 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 721 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 722 =>	"11111000",	-- #####...
--   =>	"00011000",	-- ...##...
 723 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xb5='\xb5
 724 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 725 =>	"11111000",	-- #####...
--   =>	"00011000",	-- ...##...
 726 =>	"11111000",	-- #####...
--   =>	"00011000",	-- ...##...
 727 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xb6='\xb6
 728 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 729 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 730 =>	"11110110",	-- ####.##.
--   =>	"00110110",	-- ..##.##.
 731 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xb7='\xb7
 732 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 733 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 734 =>	"11111110",	-- #######.
--   =>	"00110110",	-- ..##.##.
 735 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xb8='\xb8
 736 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 737 =>	"11111000",	-- #####...
--   =>	"00011000",	-- ...##...
 738 =>	"11111000",	-- #####...
--   =>	"00011000",	-- ...##...
 739 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xb9='\xb9
 740 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 741 =>	"11110110",	-- ####.##.
--   =>	"00000110",	-- .....##.
 742 =>	"11110110",	-- ####.##.
--   =>	"00110110",	-- ..##.##.
 743 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xba='\xba
 744 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 745 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 746 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 747 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xbb='\xbb
 748 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 749 =>	"11111110",	-- #######.
--   =>	"00000110",	-- .....##.
 750 =>	"11110110",	-- ####.##.
--   =>	"00110110",	-- ..##.##.
 751 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xbc='\xbc
 752 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 753 =>	"11110110",	-- ####.##.
--   =>	"00000110",	-- .....##.
 754 =>	"11111110",	-- #######.
--   =>	"00000000",	-- ........
 755 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xbd='\xbd
 756 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 757 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 758 =>	"11111110",	-- #######.
--   =>	"00000000",	-- ........
 759 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xbe='\xbe
 760 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 761 =>	"11111000",	-- #####...
--   =>	"00011000",	-- ...##...
 762 =>	"11111000",	-- #####...
--   =>	"00000000",	-- ........
 763 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xbf='\xbf
 764 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 765 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 766 =>	"11111000",	-- #####...
--   =>	"00011000",	-- ...##...
 767 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xc0='\xc0
 768 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 769 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 770 =>	"00011111",	-- ...#####
--   =>	"00000000",	-- ........
 771 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xc1='\xc1
 772 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 773 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 774 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 775 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xc2='\xc2
 776 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 777 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 778 =>	"11111111",	-- ########
--   =>	"00011000",	-- ...##...
 779 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xc3='\xc3
 780 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 781 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 782 =>	"00011111",	-- ...#####
--   =>	"00011000",	-- ...##...
 783 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xc4='\xc4
 784 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 785 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 786 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 787 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xc5='\xc5
 788 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 789 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 790 =>	"11111111",	-- ########
--   =>	"00011000",	-- ...##...
 791 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xc6='\xc6
 792 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 793 =>	"00011111",	-- ...#####
--   =>	"00011000",	-- ...##...
 794 =>	"00011111",	-- ...#####
--   =>	"00011000",	-- ...##...
 795 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xc7='\xc7
 796 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 797 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 798 =>	"00110111",	-- ..##.###
--   =>	"00110110",	-- ..##.##.
 799 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xc8='\xc8
 800 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 801 =>	"00110111",	-- ..##.###
--   =>	"00110000",	-- ..##....
 802 =>	"00111111",	-- ..######
--   =>	"00000000",	-- ........
 803 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xc9='\xc9
 804 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 805 =>	"00111111",	-- ..######
--   =>	"00110000",	-- ..##....
 806 =>	"00110111",	-- ..##.###
--   =>	"00110110",	-- ..##.##.
 807 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xca='\xca
 808 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 809 =>	"11110111",	-- ####.###
--   =>	"00000000",	-- ........
 810 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 811 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xcb='\xcb
 812 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 813 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 814 =>	"11110111",	-- ####.###
--   =>	"00110110",	-- ..##.##.
 815 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xcc='\xcc
 816 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 817 =>	"00110111",	-- ..##.###
--   =>	"00110000",	-- ..##....
 818 =>	"00110111",	-- ..##.###
--   =>	"00110110",	-- ..##.##.
 819 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xcd='\xcd
 820 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 821 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 822 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 823 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xce='\xce
 824 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 825 =>	"11110111",	-- ####.###
--   =>	"00000000",	-- ........
 826 =>	"11110111",	-- ####.###
--   =>	"00110110",	-- ..##.##.
 827 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xcf='\xcf
 828 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 829 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 830 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 831 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xd0='\xd0
 832 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 833 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 834 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 835 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xd1='\xd1
 836 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 837 =>	"11111111",	-- ########
--   =>	"00000000",	-- ........
 838 =>	"11111111",	-- ########
--   =>	"00011000",	-- ...##...
 839 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xd2='\xd2
 840 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 841 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 842 =>	"11111111",	-- ########
--   =>	"00110110",	-- ..##.##.
 843 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xd3='\xd3
 844 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 845 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 846 =>	"00111111",	-- ..######
--   =>	"00000000",	-- ........
 847 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xd4='\xd4
 848 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 849 =>	"00011111",	-- ...#####
--   =>	"00011000",	-- ...##...
 850 =>	"00011111",	-- ...#####
--   =>	"00000000",	-- ........
 851 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xd5='\xd5
 852 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 853 =>	"00011111",	-- ...#####
--   =>	"00011000",	-- ...##...
 854 =>	"00011111",	-- ...#####
--   =>	"00011000",	-- ...##...
 855 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xd6='\xd6
 856 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 857 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 858 =>	"00111111",	-- ..######
--   =>	"00110110",	-- ..##.##.
 859 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xd7='\xd7
 860 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 861 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.
 862 =>	"11111111",	-- ########
--   =>	"00110110",	-- ..##.##.
 863 =>	"00110110",	-- ..##.##.
--   =>	"00110110",	-- ..##.##.

-- char 0xd8='\xd8
 864 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 865 =>	"11111111",	-- ########
--   =>	"00011000",	-- ...##...
 866 =>	"11111111",	-- ########
--   =>	"00011000",	-- ...##...
 867 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xd9='\xd9
 868 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 869 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 870 =>	"11111000",	-- #####...
--   =>	"00000000",	-- ........
 871 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xda='\xda
 872 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 873 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 874 =>	"00011111",	-- ...#####
--   =>	"00011000",	-- ...##...
 875 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xdb='\xdb
 876 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 877 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 878 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 879 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########

-- char 0xdc='\xdc
 880 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 881 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 882 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 883 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########

-- char 0xdd='\xdd
 884 =>	"11110000",	-- ####....
--   =>	"11110000",	-- ####....
 885 =>	"11110000",	-- ####....
--   =>	"11110000",	-- ####....
 886 =>	"11110000",	-- ####....
--   =>	"11110000",	-- ####....
 887 =>	"11110000",	-- ####....
--   =>	"11110000",	-- ####....

-- char 0xde='\xde
 888 =>	"00001111",	-- ....####
--   =>	"00001111",	-- ....####
 889 =>	"00001111",	-- ....####
--   =>	"00001111",	-- ....####
 890 =>	"00001111",	-- ....####
--   =>	"00001111",	-- ....####
 891 =>	"00001111",	-- ....####
--   =>	"00001111",	-- ....####

-- char 0xdf='\xdf
 892 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 893 =>	"11111111",	-- ########
--   =>	"11111111",	-- ########
 894 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 895 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xe0='\xe0
 896 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 897 =>	"01110110",	-- .###.##.
--   =>	"11011100",	-- ##.###..
 898 =>	"11001000",	-- ##..#...
--   =>	"11011100",	-- ##.###..
 899 =>	"01110110",	-- .###.##.
--   =>	"00000000",	-- ........

-- char 0xe1='\xe1
 900 =>	"00000000",	-- ........
--   =>	"01111000",	-- .####...
 901 =>	"11001100",	-- ##..##..
--   =>	"11111000",	-- #####...
 902 =>	"11001100",	-- ##..##..
--   =>	"11111000",	-- #####...
 903 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......

-- char 0xe2='\xe2
 904 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 905 =>	"11001100",	-- ##..##..
--   =>	"11000000",	-- ##......
 906 =>	"11000000",	-- ##......
--   =>	"11000000",	-- ##......
 907 =>	"11000000",	-- ##......
--   =>	"00000000",	-- ........

-- char 0xe3='\xe3
 908 =>	"00000000",	-- ........
--   =>	"11111110",	-- #######.
 909 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 910 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 911 =>	"01101100",	-- .##.##..
--   =>	"00000000",	-- ........

-- char 0xe4='\xe4
 912 =>	"11111100",	-- ######..
--   =>	"11001100",	-- ##..##..
 913 =>	"01100000",	-- .##.....
--   =>	"00110000",	-- ..##....
 914 =>	"01100000",	-- .##.....
--   =>	"11001100",	-- ##..##..
 915 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0xe5='\xe5
 916 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 917 =>	"01111110",	-- .######.
--   =>	"11011000",	-- ##.##...
 918 =>	"11011000",	-- ##.##...
--   =>	"11011000",	-- ##.##...
 919 =>	"01110000",	-- .###....
--   =>	"00000000",	-- ........

-- char 0xe6='\xe6
 920 =>	"00000000",	-- ........
--   =>	"01100110",	-- .##..##.
 921 =>	"01100110",	-- .##..##.
--   =>	"01100110",	-- .##..##.
 922 =>	"01100110",	-- .##..##.
--   =>	"01111100",	-- .#####..
 923 =>	"01100000",	-- .##.....
--   =>	"11000000",	-- ##......

-- char 0xe7='\xe7
 924 =>	"00000000",	-- ........
--   =>	"01110110",	-- .###.##.
 925 =>	"11011100",	-- ##.###..
--   =>	"00011000",	-- ...##...
 926 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 927 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........

-- char 0xe8='\xe8
 928 =>	"11111100",	-- ######..
--   =>	"00110000",	-- ..##....
 929 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 930 =>	"11001100",	-- ##..##..
--   =>	"01111000",	-- .####...
 931 =>	"00110000",	-- ..##....
--   =>	"11111100",	-- ######..

-- char 0xe9='\xe9
 932 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 933 =>	"11000110",	-- ##...##.
--   =>	"11111110",	-- #######.
 934 =>	"11000110",	-- ##...##.
--   =>	"01101100",	-- .##.##..
 935 =>	"00111000",	-- ..###...
--   =>	"00000000",	-- ........

-- char 0xea='\xea
 936 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 937 =>	"11000110",	-- ##...##.
--   =>	"11000110",	-- ##...##.
 938 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
 939 =>	"11101110",	-- ###.###.
--   =>	"00000000",	-- ........

-- char 0xeb='\xeb
 940 =>	"00011100",	-- ...###..
--   =>	"00110000",	-- ..##....
 941 =>	"00011000",	-- ...##...
--   =>	"01111100",	-- .#####..
 942 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 943 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........

-- char 0xec='\xec
 944 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 945 =>	"01111110",	-- .######.
--   =>	"11011011",	-- ##.##.##
 946 =>	"11011011",	-- ##.##.##
--   =>	"01111110",	-- .######.
 947 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xed='\xed
 948 =>	"00000110",	-- .....##.
--   =>	"00001100",	-- ....##..
 949 =>	"01111110",	-- .######.
--   =>	"11011011",	-- ##.##.##
 950 =>	"11011011",	-- ##.##.##
--   =>	"01111110",	-- .######.
 951 =>	"01100000",	-- .##.....
--   =>	"11000000",	-- ##......

-- char 0xee='\xee
 952 =>	"00111000",	-- ..###...
--   =>	"01100000",	-- .##.....
 953 =>	"11000000",	-- ##......
--   =>	"11111000",	-- #####...
 954 =>	"11000000",	-- ##......
--   =>	"01100000",	-- .##.....
 955 =>	"00111000",	-- ..###...
--   =>	"00000000",	-- ........

-- char 0xef='\xef
 956 =>	"01111000",	-- .####...
--   =>	"11001100",	-- ##..##..
 957 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 958 =>	"11001100",	-- ##..##..
--   =>	"11001100",	-- ##..##..
 959 =>	"11001100",	-- ##..##..
--   =>	"00000000",	-- ........

-- char 0xf0='\xf0
 960 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 961 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 962 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 963 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xf1='\xf1
 964 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 965 =>	"11111100",	-- ######..
--   =>	"00110000",	-- ..##....
 966 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........
 967 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0xf2='\xf2
 968 =>	"01100000",	-- .##.....
--   =>	"00110000",	-- ..##....
 969 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
 970 =>	"01100000",	-- .##.....
--   =>	"00000000",	-- ........
 971 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0xf3='\xf3
 972 =>	"00011000",	-- ...##...
--   =>	"00110000",	-- ..##....
 973 =>	"01100000",	-- .##.....
--   =>	"00110000",	-- ..##....
 974 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........
 975 =>	"11111100",	-- ######..
--   =>	"00000000",	-- ........

-- char 0xf4='\xf4
 976 =>	"00001110",	-- ....###.
--   =>	"00011011",	-- ...##.##
 977 =>	"00011011",	-- ...##.##
--   =>	"00011000",	-- ...##...
 978 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 979 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...

-- char 0xf5='\xf5
 980 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 981 =>	"00011000",	-- ...##...
--   =>	"00011000",	-- ...##...
 982 =>	"00011000",	-- ...##...
--   =>	"11011000",	-- ##.##...
 983 =>	"11011000",	-- ##.##...
--   =>	"01110000",	-- .###....

-- char 0xf6='\xf6
 984 =>	"00110000",	-- ..##....
--   =>	"00110000",	-- ..##....
 985 =>	"00000000",	-- ........
--   =>	"11111100",	-- ######..
 986 =>	"00000000",	-- ........
--   =>	"00110000",	-- ..##....
 987 =>	"00110000",	-- ..##....
--   =>	"00000000",	-- ........

-- char 0xf7='\xf7
 988 =>	"00000000",	-- ........
--   =>	"01110110",	-- .###.##.
 989 =>	"11011100",	-- ##.###..
--   =>	"00000000",	-- ........
 990 =>	"01110110",	-- .###.##.
--   =>	"11011100",	-- ##.###..
 991 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xf8='\xf8
 992 =>	"00111000",	-- ..###...
--   =>	"01101100",	-- .##.##..
 993 =>	"01101100",	-- .##.##..
--   =>	"00111000",	-- ..###...
 994 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 995 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xf9='\xf9
 996 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
 997 =>	"00000000",	-- ........
--   =>	"00011000",	-- ...##...
 998 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........
 999 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xfa='\xfa
1000 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1001 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1002 =>	"00011000",	-- ...##...
--   =>	"00000000",	-- ........
1003 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xfb='\xfb
1004 =>	"00001111",	-- ....####
--   =>	"00001100",	-- ....##..
1005 =>	"00001100",	-- ....##..
--   =>	"00001100",	-- ....##..
1006 =>	"11101100",	-- ###.##..
--   =>	"01101100",	-- .##.##..
1007 =>	"00111100",	-- ..####..
--   =>	"00011100",	-- ...###..

-- char 0xfc='\xfc
1008 =>	"01111000",	-- .####...
--   =>	"01101100",	-- .##.##..
1009 =>	"01101100",	-- .##.##..
--   =>	"01101100",	-- .##.##..
1010 =>	"01101100",	-- .##.##..
--   =>	"00000000",	-- ........
1011 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xfd='\xfd
1012 =>	"01110000",	-- .###....
--   =>	"00011000",	-- ...##...
1013 =>	"00110000",	-- ..##....
--   =>	"01100000",	-- .##.....
1014 =>	"01111000",	-- .####...
--   =>	"00000000",	-- ........
1015 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xfe='\xfe
1016 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1017 =>	"00111100",	-- ..####..
--   =>	"00111100",	-- ..####..
1018 =>	"00111100",	-- ..####..
--   =>	"00111100",	-- ..####..
1019 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........

-- char 0xff='\xff
1020 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1021 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1022 =>	"00000000",	-- ........
--   =>	"00000000",	-- ........
1023 =>	"00000000"	-- ........
--   =>	"00000000",	-- ........
);
	attribute syn_ramstyle: string;
	attribute syn_ramstyle of mem: signal is "no_rw_check";
begin
	process (clka_i) -- Using port a.
	begin
	if (rising_edge(clka_i)) then
		if (wea_i = '1') then
		mem(conv_integer(addra_i)) <= dina_i;
			-- Using address bus a.
		end if;
		douta_o <= mem(conv_integer(addra_i));
	end if;
	end process;
	process (clkb_i) -- Using port b.
	begin
	if (rising_edge(clkb_i)) then
		if (web_i = '1') then
		mem(conv_integer(addrb_i)) <= dinb_i;
			-- Using address bus b.
		end if;
		doutb_o <= mem(conv_integer(addrb_i));
	end if;
	end process;
end rtl;
