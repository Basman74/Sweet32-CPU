library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
  
entity Sweet32_SRAM_lower is

   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      addr_i  : in  std_logic_vector(12 downto 0);
      write_i : in  std_logic_vector(7 downto 0);
      read_o  : out std_logic_vector(7 downto 0)
	);
end entity Sweet32_SRAM_lower;

architecture behavioral of Sweet32_SRAM_lower is
   type ram_type is array(8191 downto 0) of std_logic_vector(7 downto 0);
   signal addr_r  : std_logic_vector(12 downto 0);

   signal ram : ram_type :=
(
 
 -- Test program, lower byte (LSB) of 16-bit (byte-addressable) ROM

   0 => x"D0",
   1 => x"03",
   2 => x"00",
   3 => x"00",
   4 => x"E0",
   5 => x"7C",
   6 => x"ED",
   7 => x"1E",
   8 => x"E4",
   9 => x"1E",
  10 => x"E4",
  11 => x"1E",
  12 => x"E4",
  13 => x"1E",
  14 => x"E4",
  15 => x"1E",
  16 => x"E4",
  17 => x"1E",
  18 => x"E4",
  19 => x"1E",
  20 => x"E4",
  21 => x"1E",
  22 => x"E4",
  23 => x"1E",
  24 => x"E4",
  25 => x"1E",
  26 => x"E4",
  27 => x"1E",
  28 => x"E4",
  29 => x"1E",
  30 => x"E4",
  31 => x"1E",
  32 => x"E4",
  33 => x"1E",
  34 => x"E4",
  35 => x"00",
  36 => x"40",
  37 => x"0D",
  38 => x"1E",
  39 => x"E4",
  40 => x"1E",
  41 => x"E0",
  42 => x"C0",
  43 => x"00",
  44 => x"00",
  45 => x"00",
  46 => x"10",
  47 => x"08",
  48 => x"01",
  49 => x"31",
  50 => x"30",
  51 => x"6F",
  52 => x"60",
  53 => x"BC",
  54 => x"6D",
  55 => x"46",
  56 => x"50",
  57 => x"79",
  58 => x"F2",
  59 => x"E5",
  60 => x"00",
  61 => x"10",
  62 => x"00",
  63 => x"01",
  64 => x"E0",
  65 => x"40",
  66 => x"ED",
  67 => x"F0",
  68 => x"7C",
  69 => x"FD",
  70 => x"D6",
  71 => x"0F",
  72 => x"F4",
  73 => x"1F",
  74 => x"F4",
  75 => x"2F",
  76 => x"F4",
  77 => x"3F",
  78 => x"F4",
  79 => x"4F",
  80 => x"F4",
  81 => x"5F",
  82 => x"F4",
  83 => x"6F",
  84 => x"F4",
  85 => x"7F",
  86 => x"F4",
  87 => x"8F",
  88 => x"F4",
  89 => x"9F",
  90 => x"F4",
  91 => x"AF",
  92 => x"F4",
  93 => x"BF",
  94 => x"F4",
  95 => x"CF",
  96 => x"F0",
  97 => x"0D",
  98 => x"10",
  99 => x"40",
 100 => x"1D",
 101 => x"0F",
 102 => x"10",
 103 => x"00",
 104 => x"10",
 105 => x"00",
 106 => x"BC",
 107 => x"0D",
 108 => x"10",
 109 => x"00",
 110 => x"78",
 111 => x"0D",
 112 => x"10",
 113 => x"30",
 114 => x"E4",
 115 => x"F2",
 116 => x"C8",
 117 => x"50",
 118 => x"60",
 119 => x"76",
 120 => x"7D",
 121 => x"77",
 122 => x"66",
 123 => x"6F",
 124 => x"30",
 125 => x"FF",
 126 => x"45",
 127 => x"52",
 128 => x"F2",
 129 => x"DE",
 130 => x"30",
 131 => x"6F",
 132 => x"46",
 133 => x"F9",
 134 => x"07",
 135 => x"00",
 136 => x"0D",
 137 => x"F2",
 138 => x"73",
 139 => x"3F",
 140 => x"F2",
 141 => x"C0",
 142 => x"30",
 143 => x"F2",
 144 => x"6D",
 145 => x"30",
 146 => x"17",
 147 => x"F2",
 148 => x"A8",
 149 => x"30",
 150 => x"08",
 151 => x"F2",
 152 => x"A4",
 153 => x"F2",
 154 => x"C3",
 155 => x"FA",
 156 => x"02",
 157 => x"00",
 158 => x"00",
 159 => x"21",
 160 => x"04",
 161 => x"00",
 162 => x"00",
 163 => x"20",
 164 => x"0D",
 165 => x"00",
 166 => x"00",
 167 => x"53",
 168 => x"07",
 169 => x"00",
 170 => x"00",
 171 => x"49",
 172 => x"05",
 173 => x"00",
 174 => x"00",
 175 => x"59",
 176 => x"02",
 177 => x"00",
 178 => x"00",
 179 => x"17",
 180 => x"0C",
 181 => x"00",
 182 => x"00",
 183 => x"6D",
 184 => x"08",
 185 => x"00",
 186 => x"00",
 187 => x"9B",
 188 => x"0D",
 189 => x"00",
 190 => x"00",
 191 => x"15",
 192 => x"30",
 193 => x"0C",
 194 => x"7A",
 195 => x"EC",
 196 => x"1E",
 197 => x"30",
 198 => x"91",
 199 => x"F2",
 200 => x"74",
 201 => x"90",
 202 => x"78",
 203 => x"9D",
 204 => x"39",
 205 => x"48",
 206 => x"F2",
 207 => x"B7",
 208 => x"C0",
 209 => x"26",
 210 => x"60",
 211 => x"07",
 212 => x"EC",
 213 => x"1E",
 214 => x"90",
 215 => x"78",
 216 => x"9D",
 217 => x"69",
 218 => x"00",
 219 => x"70",
 220 => x"80",
 221 => x"30",
 222 => x"99",
 223 => x"40",
 224 => x"50",
 225 => x"82",
 226 => x"F2",
 227 => x"3D",
 228 => x"36",
 229 => x"61",
 230 => x"81",
 231 => x"F2",
 232 => x"1D",
 233 => x"07",
 234 => x"00",
 235 => x"08",
 236 => x"30",
 237 => x"F2",
 238 => x"5F",
 239 => x"0F",
 240 => x"40",
 241 => x"F3",
 242 => x"EB",
 243 => x"90",
 244 => x"78",
 245 => x"9D",
 246 => x"19",
 247 => x"FE",
 248 => x"E4",
 249 => x"0F",
 250 => x"EC",
 251 => x"1E",
 252 => x"30",
 253 => x"A1",
 254 => x"F2",
 255 => x"3D",
 256 => x"90",
 257 => x"78",
 258 => x"9D",
 259 => x"39",
 260 => x"48",
 261 => x"F2",
 262 => x"80",
 263 => x"C0",
 264 => x"19",
 265 => x"60",
 266 => x"30",
 267 => x"99",
 268 => x"40",
 269 => x"50",
 270 => x"82",
 271 => x"F2",
 272 => x"10",
 273 => x"36",
 274 => x"F2",
 275 => x"F2",
 276 => x"3D",
 277 => x"F2",
 278 => x"37",
 279 => x"36",
 280 => x"42",
 281 => x"F2",
 282 => x"6C",
 283 => x"C0",
 284 => x"05",
 285 => x"26",
 286 => x"61",
 287 => x"19",
 288 => x"EA",
 289 => x"FE",
 290 => x"E4",
 291 => x"0F",
 292 => x"EC",
 293 => x"1E",
 294 => x"30",
 295 => x"D0",
 296 => x"F2",
 297 => x"13",
 298 => x"90",
 299 => x"78",
 300 => x"9D",
 301 => x"39",
 302 => x"48",
 303 => x"F2",
 304 => x"56",
 305 => x"C0",
 306 => x"8B",
 307 => x"60",
 308 => x"07",
 309 => x"EC",
 310 => x"1E",
 311 => x"90",
 312 => x"78",
 313 => x"9D",
 314 => x"69",
 315 => x"0C",
 316 => x"70",
 317 => x"30",
 318 => x"99",
 319 => x"40",
 320 => x"50",
 321 => x"82",
 322 => x"F2",
 323 => x"DD",
 324 => x"80",
 325 => x"AE",
 326 => x"8D",
 327 => x"36",
 328 => x"08",
 329 => x"30",
 330 => x"82",
 331 => x"08",
 332 => x"03",
 333 => x"00",
 334 => x"04",
 335 => x"84",
 336 => x"86",
 337 => x"F6",
 338 => x"36",
 339 => x"F2",
 340 => x"A9",
 341 => x"30",
 342 => x"F2",
 343 => x"F6",
 344 => x"83",
 345 => x"48",
 346 => x"C1",
 347 => x"05",
 348 => x"30",
 349 => x"90",
 350 => x"F1",
 351 => x"DD",
 352 => x"32",
 353 => x"33",
 354 => x"F2",
 355 => x"9A",
 356 => x"48",
 357 => x"C0",
 358 => x"05",
 359 => x"30",
 360 => x"94",
 361 => x"F6",
 362 => x"D2",
 363 => x"34",
 364 => x"33",
 365 => x"F2",
 366 => x"8F",
 367 => x"30",
 368 => x"F2",
 369 => x"DC",
 370 => x"81",
 371 => x"30",
 372 => x"46",
 373 => x"F2",
 374 => x"B9",
 375 => x"30",
 376 => x"96",
 377 => x"F2",
 378 => x"C2",
 379 => x"8E",
 380 => x"28",
 381 => x"36",
 382 => x"40",
 383 => x"11",
 384 => x"22",
 385 => x"02",
 386 => x"31",
 387 => x"22",
 388 => x"06",
 389 => x"0F",
 390 => x"30",
 391 => x"F2",
 392 => x"B1",
 393 => x"2A",
 394 => x"22",
 395 => x"0A",
 396 => x"00",
 397 => x"30",
 398 => x"33",
 399 => x"33",
 400 => x"33",
 401 => x"33",
 402 => x"F2",
 403 => x"A6",
 404 => x"1F",
 405 => x"22",
 406 => x"0D",
 407 => x"00",
 408 => x"FF",
 409 => x"30",
 410 => x"8B",
 411 => x"03",
 412 => x"00",
 413 => x"30",
 414 => x"33",
 415 => x"34",
 416 => x"F2",
 417 => x"54",
 418 => x"11",
 419 => x"22",
 420 => x"14",
 421 => x"00",
 422 => x"FF",
 423 => x"30",
 424 => x"33",
 425 => x"12",
 426 => x"11",
 427 => x"31",
 428 => x"9B",
 429 => x"05",
 430 => x"00",
 431 => x"00",
 432 => x"00",
 433 => x"30",
 434 => x"33",
 435 => x"34",
 436 => x"32",
 437 => x"F2",
 438 => x"3F",
 439 => x"FC",
 440 => x"22",
 441 => x"10",
 442 => x"36",
 443 => x"0F",
 444 => x"30",
 445 => x"F2",
 446 => x"7B",
 447 => x"3C",
 448 => x"F2",
 449 => x"8C",
 450 => x"36",
 451 => x"0F",
 452 => x"33",
 453 => x"30",
 454 => x"F2",
 455 => x"72",
 456 => x"EB",
 457 => x"22",
 458 => x"10",
 459 => x"0F",
 460 => x"33",
 461 => x"30",
 462 => x"F2",
 463 => x"6A",
 464 => x"30",
 465 => x"7F",
 466 => x"F2",
 467 => x"69",
 468 => x"36",
 469 => x"0F",
 470 => x"30",
 471 => x"F2",
 472 => x"2D",
 473 => x"DA",
 474 => x"22",
 475 => x"09",
 476 => x"00",
 477 => x"30",
 478 => x"33",
 479 => x"33",
 480 => x"33",
 481 => x"33",
 482 => x"FD",
 483 => x"56",
 484 => x"22",
 485 => x"12",
 486 => x"00",
 487 => x"30",
 488 => x"33",
 489 => x"33",
 490 => x"33",
 491 => x"33",
 492 => x"F2",
 493 => x"4C",
 494 => x"3C",
 495 => x"F2",
 496 => x"5D",
 497 => x"36",
 498 => x"0F",
 499 => x"30",
 500 => x"F2",
 501 => x"44",
 502 => x"BD",
 503 => x"22",
 504 => x"0F",
 505 => x"00",
 506 => x"30",
 507 => x"33",
 508 => x"33",
 509 => x"33",
 510 => x"33",
 511 => x"F2",
 512 => x"39",
 513 => x"3C",
 514 => x"F2",
 515 => x"4A",
 516 => x"30",
 517 => x"FC",
 518 => x"47",
 519 => x"22",
 520 => x"04",
 521 => x"30",
 522 => x"F0",
 523 => x"42",
 524 => x"22",
 525 => x"1B",
 526 => x"00",
 527 => x"30",
 528 => x"33",
 529 => x"33",
 530 => x"33",
 531 => x"33",
 532 => x"F2",
 533 => x"24",
 534 => x"30",
 535 => x"7F",
 536 => x"F2",
 537 => x"23",
 538 => x"16",
 539 => x"0F",
 540 => x"30",
 541 => x"00",
 542 => x"00",
 543 => x"10",
 544 => x"11",
 545 => x"11",
 546 => x"11",
 547 => x"11",
 548 => x"31",
 549 => x"F2",
 550 => x"DF",
 551 => x"8C",
 552 => x"22",
 553 => x"20",
 554 => x"00",
 555 => x"30",
 556 => x"33",
 557 => x"33",
 558 => x"33",
 559 => x"33",
 560 => x"F2",
 561 => x"08",
 562 => x"3C",
 563 => x"F2",
 564 => x"19",
 565 => x"16",
 566 => x"0F",
 567 => x"30",
 568 => x"00",
 569 => x"00",
 570 => x"10",
 571 => x"11",
 572 => x"11",
 573 => x"11",
 574 => x"11",
 575 => x"31",
 576 => x"87",
 577 => x"04",
 578 => x"0F",
 579 => x"00",
 580 => x"30",
 581 => x"33",
 582 => x"36",
 583 => x"FC",
 584 => x"AD",
 585 => x"22",
 586 => x"11",
 587 => x"00",
 588 => x"30",
 589 => x"33",
 590 => x"33",
 591 => x"33",
 592 => x"33",
 593 => x"F2",
 594 => x"E7",
 595 => x"30",
 596 => x"7F",
 597 => x"F2",
 598 => x"E6",
 599 => x"32",
 600 => x"33",
 601 => x"FA",
 602 => x"A3",
 603 => x"22",
 604 => x"11",
 605 => x"00",
 606 => x"30",
 607 => x"33",
 608 => x"33",
 609 => x"33",
 610 => x"33",
 611 => x"F2",
 612 => x"D5",
 613 => x"30",
 614 => x"7F",
 615 => x"F2",
 616 => x"D4",
 617 => x"32",
 618 => x"33",
 619 => x"F8",
 620 => x"89",
 621 => x"22",
 622 => x"13",
 623 => x"00",
 624 => x"30",
 625 => x"33",
 626 => x"33",
 627 => x"33",
 628 => x"33",
 629 => x"F2",
 630 => x"C3",
 631 => x"3C",
 632 => x"F2",
 633 => x"D4",
 634 => x"36",
 635 => x"0F",
 636 => x"33",
 637 => x"30",
 638 => x"F2",
 639 => x"BA",
 640 => x"6E",
 641 => x"22",
 642 => x"0D",
 643 => x"00",
 644 => x"30",
 645 => x"33",
 646 => x"33",
 647 => x"33",
 648 => x"33",
 649 => x"F2",
 650 => x"AF",
 651 => x"3C",
 652 => x"F2",
 653 => x"C0",
 654 => x"2C",
 655 => x"00",
 656 => x"30",
 657 => x"33",
 658 => x"33",
 659 => x"33",
 660 => x"33",
 661 => x"F2",
 662 => x"A3",
 663 => x"3C",
 664 => x"F2",
 665 => x"B4",
 666 => x"36",
 667 => x"0F",
 668 => x"33",
 669 => x"30",
 670 => x"F2",
 671 => x"9A",
 672 => x"30",
 673 => x"7F",
 674 => x"F2",
 675 => x"99",
 676 => x"36",
 677 => x"0F",
 678 => x"30",
 679 => x"83",
 680 => x"09",
 681 => x"50",
 682 => x"3D",
 683 => x"F2",
 684 => x"A1",
 685 => x"07",
 686 => x"35",
 687 => x"30",
 688 => x"31",
 689 => x"F2",
 690 => x"62",
 691 => x"81",
 692 => x"08",
 693 => x"00",
 694 => x"60",
 695 => x"07",
 696 => x"85",
 697 => x"90",
 698 => x"78",
 699 => x"9D",
 700 => x"19",
 701 => x"FE",
 702 => x"E4",
 703 => x"0F",
 704 => x"EC",
 705 => x"1E",
 706 => x"04",
 707 => x"60",
 708 => x"30",
 709 => x"97",
 710 => x"F2",
 711 => x"75",
 712 => x"80",
 713 => x"30",
 714 => x"21",
 715 => x"F2",
 716 => x"70",
 717 => x"30",
 718 => x"F2",
 719 => x"2E",
 720 => x"F2",
 721 => x"7B",
 722 => x"F2",
 723 => x"8A",
 724 => x"50",
 725 => x"16",
 726 => x"61",
 727 => x"CF",
 728 => x"F1",
 729 => x"04",
 730 => x"00",
 731 => x"30",
 732 => x"F2",
 733 => x"70",
 734 => x"30",
 735 => x"F2",
 736 => x"6D",
 737 => x"05",
 738 => x"00",
 739 => x"40",
 740 => x"E5",
 741 => x"81",
 742 => x"81",
 743 => x"E2",
 744 => x"30",
 745 => x"5F",
 746 => x"F2",
 747 => x"51",
 748 => x"30",
 749 => x"F2",
 750 => x"0F",
 751 => x"F2",
 752 => x"5C",
 753 => x"FE",
 754 => x"E4",
 755 => x"0F",
 756 => x"EC",
 757 => x"1E",
 758 => x"30",
 759 => x"9D",
 760 => x"F4",
 761 => x"43",
 762 => x"50",
 763 => x"BC",
 764 => x"5D",
 765 => x"35",
 766 => x"48",
 767 => x"F2",
 768 => x"86",
 769 => x"C0",
 770 => x"03",
 771 => x"15",
 772 => x"2E",
 773 => x"FE",
 774 => x"E4",
 775 => x"0F",
 776 => x"EC",
 777 => x"1E",
 778 => x"34",
 779 => x"33",
 780 => x"41",
 781 => x"0C",
 782 => x"C9",
 783 => x"07",
 784 => x"33",
 785 => x"FC",
 786 => x"30",
 787 => x"D6",
 788 => x"F2",
 789 => x"27",
 790 => x"B0",
 791 => x"50",
 792 => x"F2",
 793 => x"51",
 794 => x"05",
 795 => x"02",
 796 => x"40",
 797 => x"03",
 798 => x"B1",
 799 => x"F9",
 800 => x"03",
 801 => x"02",
 802 => x"00",
 803 => x"0A",
 804 => x"0B",
 805 => x"02",
 806 => x"00",
 807 => x"83",
 808 => x"51",
 809 => x"B0",
 810 => x"82",
 811 => x"ED",
 812 => x"3C",
 813 => x"F2",
 814 => x"3C",
 815 => x"07",
 816 => x"02",
 817 => x"40",
 818 => x"36",
 819 => x"F2",
 820 => x"7E",
 821 => x"00",
 822 => x"33",
 823 => x"02",
 824 => x"40",
 825 => x"2F",
 826 => x"F2",
 827 => x"77",
 828 => x"00",
 829 => x"76",
 830 => x"02",
 831 => x"40",
 832 => x"28",
 833 => x"80",
 834 => x"BC",
 835 => x"8D",
 836 => x"F2",
 837 => x"79",
 838 => x"3D",
 839 => x"0C",
 840 => x"88",
 841 => x"FE",
 842 => x"0C",
 843 => x"46",
 844 => x"18",
 845 => x"06",
 846 => x"68",
 847 => x"F2",
 848 => x"6E",
 849 => x"00",
 850 => x"FF",
 851 => x"FF",
 852 => x"06",
 853 => x"13",
 854 => x"3A",
 855 => x"0C",
 856 => x"88",
 857 => x"FE",
 858 => x"0C",
 859 => x"70",
 860 => x"88",
 861 => x"F2",
 862 => x"54",
 863 => x"40",
 864 => x"08",
 865 => x"82",
 866 => x"7F",
 867 => x"07",
 868 => x"09",
 869 => x"3E",
 870 => x"F7",
 871 => x"E6",
 872 => x"B0",
 873 => x"30",
 874 => x"01",
 875 => x"FF",
 876 => x"D0",
 877 => x"F2",
 878 => x"44",
 879 => x"00",
 880 => x"4E",
 881 => x"02",
 882 => x"40",
 883 => x"F5",
 884 => x"F2",
 885 => x"3D",
 886 => x"70",
 887 => x"30",
 888 => x"F2",
 889 => x"40",
 890 => x"BC",
 891 => x"4D",
 892 => x"44",
 893 => x"50",
 894 => x"F2",
 895 => x"A1",
 896 => x"3D",
 897 => x"F2",
 898 => x"CB",
 899 => x"40",
 900 => x"BC",
 901 => x"4D",
 902 => x"44",
 903 => x"34",
 904 => x"F2",
 905 => x"6C",
 906 => x"30",
 907 => x"FB",
 908 => x"F2",
 909 => x"AF",
 910 => x"00",
 911 => x"BC",
 912 => x"0D",
 913 => x"50",
 914 => x"30",
 915 => x"FF",
 916 => x"45",
 917 => x"52",
 918 => x"F2",
 919 => x"C8",
 920 => x"30",
 921 => x"6F",
 922 => x"46",
 923 => x"F9",
 924 => x"80",
 925 => x"30",
 926 => x"F2",
 927 => x"5E",
 928 => x"30",
 929 => x"13",
 930 => x"F8",
 931 => x"07",
 932 => x"00",
 933 => x"04",
 934 => x"30",
 935 => x"17",
 936 => x"F0",
 937 => x"93",
 938 => x"BF",
 939 => x"0B",
 940 => x"86",
 941 => x"F2",
 942 => x"9E",
 943 => x"FE",
 944 => x"E4",
 945 => x"0F",
 946 => x"EC",
 947 => x"1E",
 948 => x"F2",
 949 => x"B5",
 950 => x"10",
 951 => x"F2",
 952 => x"B2",
 953 => x"22",
 954 => x"21",
 955 => x"FE",
 956 => x"E4",
 957 => x"0F",
 958 => x"EC",
 959 => x"1E",
 960 => x"F2",
 961 => x"F1",
 962 => x"60",
 963 => x"F2",
 964 => x"EE",
 965 => x"22",
 966 => x"62",
 967 => x"FE",
 968 => x"E4",
 969 => x"0F",
 970 => x"EC",
 971 => x"1E",
 972 => x"30",
 973 => x"A9",
 974 => x"F2",
 975 => x"6D",
 976 => x"60",
 977 => x"30",
 978 => x"09",
 979 => x"F3",
 980 => x"00",
 981 => x"78",
 982 => x"30",
 983 => x"F2",
 984 => x"57",
 985 => x"50",
 986 => x"7C",
 987 => x"5D",
 988 => x"06",
 989 => x"00",
 990 => x"50",
 991 => x"35",
 992 => x"F2",
 993 => x"14",
 994 => x"64",
 995 => x"F7",
 996 => x"00",
 997 => x"06",
 998 => x"66",
 999 => x"30",
1000 => x"F9",
1001 => x"64",
1002 => x"61",
1003 => x"0F",
1004 => x"60",
1005 => x"03",
1006 => x"40",
1007 => x"E2",
1008 => x"30",
1009 => x"ED",
1010 => x"F2",
1011 => x"49",
1012 => x"00",
1013 => x"BC",
1014 => x"0D",
1015 => x"30",
1016 => x"F2",
1017 => x"FC",
1018 => x"F2",
1019 => x"51",
1020 => x"30",
1021 => x"B4",
1022 => x"F2",
1023 => x"3D",
1024 => x"3C",
1025 => x"42",
1026 => x"F2",
1027 => x"83",
1028 => x"C0",
1029 => x"27",
1030 => x"70",
1031 => x"0C",
1032 => x"00",
1033 => x"00",
1034 => x"76",
1035 => x"00",
1036 => x"16",
1037 => x"07",
1038 => x"77",
1039 => x"00",
1040 => x"01",
1041 => x"07",
1042 => x"1A",
1043 => x"30",
1044 => x"89",
1045 => x"F2",
1046 => x"26",
1047 => x"30",
1048 => x"09",
1049 => x"F3",
1050 => x"00",
1051 => x"32",
1052 => x"30",
1053 => x"F2",
1054 => x"11",
1055 => x"10",
1056 => x"7C",
1057 => x"1D",
1058 => x"07",
1059 => x"00",
1060 => x"70",
1061 => x"37",
1062 => x"48",
1063 => x"F2",
1064 => x"5E",
1065 => x"C0",
1066 => x"02",
1067 => x"17",
1068 => x"FE",
1069 => x"E4",
1070 => x"0F",
1071 => x"EC",
1072 => x"1E",
1073 => x"FF",
1074 => x"07",
1075 => x"3D",
1076 => x"FF",
1077 => x"18",
1078 => x"FE",
1079 => x"E4",
1080 => x"0F",
1081 => x"EC",
1082 => x"1E",
1083 => x"40",
1084 => x"00",
1085 => x"00",
1086 => x"40",
1087 => x"05",
1088 => x"30",
1089 => x"ED",
1090 => x"F1",
1091 => x"F9",
1092 => x"32",
1093 => x"F2",
1094 => x"07",
1095 => x"31",
1096 => x"0A",
1097 => x"F3",
1098 => x"04",
1099 => x"02",
1100 => x"30",
1101 => x"0A",
1102 => x"14",
1103 => x"33",
1104 => x"00",
1105 => x"F2",
1106 => x"C2",
1107 => x"FE",
1108 => x"E4",
1109 => x"0F",
1110 => x"EC",
1111 => x"1E",
1112 => x"30",
1113 => x"9B",
1114 => x"F2",
1115 => x"E1",
1116 => x"FE",
1117 => x"E4",
1118 => x"0F",
1119 => x"EC",
1120 => x"1E",
1121 => x"EC",
1122 => x"1E",
1123 => x"54",
1124 => x"0F",
1125 => x"40",
1126 => x"F2",
1127 => x"08",
1128 => x"30",
1129 => x"0F",
1130 => x"40",
1131 => x"5E",
1132 => x"E4",
1133 => x"FE",
1134 => x"E4",
1135 => x"13",
1136 => x"0F",
1137 => x"10",
1138 => x"41",
1139 => x"14",
1140 => x"11",
1141 => x"11",
1142 => x"11",
1143 => x"41",
1144 => x"23",
1145 => x"00",
1146 => x"20",
1147 => x"24",
1148 => x"00",
1149 => x"40",
1150 => x"24",
1151 => x"00",
1152 => x"40",
1153 => x"24",
1154 => x"00",
1155 => x"FF",
1156 => x"20",
1157 => x"0F",
1158 => x"EC",
1159 => x"1E",
1160 => x"EC",
1161 => x"1E",
1162 => x"EC",
1163 => x"1E",
1164 => x"EC",
1165 => x"1E",
1166 => x"EC",
1167 => x"1E",
1168 => x"EC",
1169 => x"1E",
1170 => x"50",
1171 => x"60",
1172 => x"70",
1173 => x"80",
1174 => x"40",
1175 => x"90",
1176 => x"F2",
1177 => x"C4",
1178 => x"0B",
1179 => x"00",
1180 => x"00",
1181 => x"30",
1182 => x"0D",
1183 => x"00",
1184 => x"00",
1185 => x"30",
1186 => x"08",
1187 => x"00",
1188 => x"00",
1189 => x"1D",
1190 => x"09",
1191 => x"00",
1192 => x"00",
1193 => x"26",
1194 => x"30",
1195 => x"00",
1196 => x"22",
1197 => x"00",
1198 => x"0A",
1199 => x"17",
1200 => x"02",
1201 => x"22",
1202 => x"00",
1203 => x"0F",
1204 => x"00",
1205 => x"40",
1206 => x"E1",
1207 => x"07",
1208 => x"00",
1209 => x"DE",
1210 => x"71",
1211 => x"55",
1212 => x"55",
1213 => x"55",
1214 => x"55",
1215 => x"52",
1216 => x"F7",
1217 => x"8C",
1218 => x"07",
1219 => x"D4",
1220 => x"55",
1221 => x"55",
1222 => x"55",
1223 => x"55",
1224 => x"7F",
1225 => x"30",
1226 => x"85",
1227 => x"FC",
1228 => x"70",
1229 => x"41",
1230 => x"05",
1231 => x"91",
1232 => x"50",
1233 => x"07",
1234 => x"50",
1235 => x"07",
1236 => x"06",
1237 => x"7F",
1238 => x"30",
1239 => x"85",
1240 => x"FB",
1241 => x"63",
1242 => x"44",
1243 => x"0A",
1244 => x"70",
1245 => x"30",
1246 => x"F7",
1247 => x"83",
1248 => x"02",
1249 => x"14",
1250 => x"C2",
1251 => x"1A",
1252 => x"21",
1253 => x"49",
1254 => x"B1",
1255 => x"20",
1256 => x"5E",
1257 => x"E4",
1258 => x"6E",
1259 => x"E4",
1260 => x"7E",
1261 => x"E4",
1262 => x"8E",
1263 => x"E4",
1264 => x"9E",
1265 => x"E4",
1266 => x"FE",
1267 => x"E4",
1268 => x"0F",
1269 => x"EC",
1270 => x"1E",
1271 => x"33",
1272 => x"F2",
1273 => x"04",
1274 => x"33",
1275 => x"FE",
1276 => x"E4",
1277 => x"EC",
1278 => x"1E",
1279 => x"33",
1280 => x"F2",
1281 => x"04",
1282 => x"33",
1283 => x"FE",
1284 => x"E4",
1285 => x"13",
1286 => x"11",
1287 => x"11",
1288 => x"11",
1289 => x"0F",
1290 => x"10",
1291 => x"00",
1292 => x"10",
1293 => x"0A",
1294 => x"01",
1295 => x"17",
1296 => x"0C",
1297 => x"88",
1298 => x"FE",
1299 => x"0C",
1300 => x"0F",
1301 => x"10",
1302 => x"00",
1303 => x"10",
1304 => x"0A",
1305 => x"01",
1306 => x"17",
1307 => x"0C",
1308 => x"88",
1309 => x"FE",
1310 => x"0C",
1311 => x"0F",
1312 => x"EC",
1313 => x"1E",
1314 => x"F2",
1315 => x"19",
1316 => x"30",
1317 => x"F2",
1318 => x"CF",
1319 => x"30",
1320 => x"03",
1321 => x"03",
1322 => x"F2",
1323 => x"11",
1324 => x"FE",
1325 => x"E4",
1326 => x"0F",
1327 => x"EC",
1328 => x"1E",
1329 => x"20",
1330 => x"32",
1331 => x"F2",
1332 => x"19",
1333 => x"21",
1334 => x"4F",
1335 => x"44",
1336 => x"FA",
1337 => x"FE",
1338 => x"E4",
1339 => x"0F",
1340 => x"EC",
1341 => x"1E",
1342 => x"EC",
1343 => x"1E",
1344 => x"2D",
1345 => x"32",
1346 => x"21",
1347 => x"03",
1348 => x"03",
1349 => x"FC",
1350 => x"07",
1351 => x"4E",
1352 => x"E4",
1353 => x"FE",
1354 => x"E4",
1355 => x"0F",
1356 => x"3A",
1357 => x"0F",
1358 => x"30",
1359 => x"0A",
1360 => x"03",
1361 => x"40",
1362 => x"06",
1363 => x"0C",
1364 => x"88",
1365 => x"FE",
1366 => x"0D",
1367 => x"0C",
1368 => x"0C",
1369 => x"88",
1370 => x"FE",
1371 => x"0C",
1372 => x"0F",
1373 => x"EC",
1374 => x"1E",
1375 => x"F2",
1376 => x"0A",
1377 => x"00",
1378 => x"00",
1379 => x"04",
1380 => x"00",
1381 => x"22",
1382 => x"00",
1383 => x"FE",
1384 => x"E4",
1385 => x"0F",
1386 => x"2C",
1387 => x"89",
1388 => x"FE",
1389 => x"02",
1390 => x"00",
1391 => x"0F",
1392 => x"20",
1393 => x"0F",
1394 => x"0A",
1395 => x"77",
1396 => x"65",
1397 => x"33",
1398 => x"20",
1399 => x"6F",
1400 => x"69",
1401 => x"6F",
1402 => x"2F",
1403 => x"6F",
1404 => x"64",
1405 => x"72",
1406 => x"76",
1407 => x"2E",
1408 => x"32",
1409 => x"62",
1410 => x"74",
1411 => x"0A",
1412 => x"0A",
1413 => x"20",
1414 => x"3F",
1415 => x"0A",
1416 => x"44",
1417 => x"2D",
1418 => x"44",
1419 => x"6D",
1420 => x"20",
1421 => x"65",
1422 => x"6F",
1423 => x"79",
1424 => x"20",
1425 => x"20",
1426 => x"20",
1427 => x"6F",
1428 => x"69",
1429 => x"79",
1430 => x"6D",
1431 => x"6D",
1432 => x"72",
1433 => x"0A",
1434 => x"47",
1435 => x"2D",
1436 => x"47",
1437 => x"20",
1438 => x"65",
1439 => x"65",
1440 => x"75",
1441 => x"65",
1442 => x"0A",
1443 => x"52",
1444 => x"2D",
1445 => x"52",
1446 => x"67",
1447 => x"73",
1448 => x"65",
1449 => x"73",
1450 => x"20",
1451 => x"20",
1452 => x"20",
1453 => x"61",
1454 => x"64",
1455 => x"72",
1456 => x"74",
1457 => x"20",
1458 => x"65",
1459 => x"0A",
1460 => x"55",
1461 => x"2D",
1462 => x"55",
1463 => x"6C",
1464 => x"61",
1465 => x"20",
1466 => x"57",
1467 => x"20",
1468 => x"69",
1469 => x"65",
1470 => x"28",
1471 => x"72",
1472 => x"73",
1473 => x"6E",
1474 => x"20",
1475 => x"74",
1476 => x"70",
1477 => x"6F",
1478 => x"70",
1479 => x"29",
1480 => x"00",
1481 => x"75",
1482 => x"70",
1483 => x"00",
1484 => x"61",
1485 => x"64",
1486 => x"00",
1487 => x"6F",
1488 => x"00",
1489 => x"6F",
1490 => x"69",
1491 => x"79",
1492 => x"00",
1493 => x"65",
1494 => x"69",
1495 => x"74",
1496 => x"72",
1497 => x"0A",
1498 => x"4D",
1499 => x"64",
1500 => x"66",
1501 => x"20",
1502 => x"65",
1503 => x"20",
1504 => x"2D",
1505 => x"35",
1506 => x"28",
1507 => x"20",
1508 => x"6F",
1509 => x"20",
1510 => x"63",
1511 => x"20",
1512 => x"4C",
1513 => x"73",
1514 => x"20",
1515 => x"55",
1516 => x"6C",
1517 => x"61",
1518 => x"0A",
1519 => x"77",
1520 => x"69",
1521 => x"69",
1522 => x"67",
1523 => x"53",
1524 => x"45",
1525 => x"2E",
1526 => x"00",
1527 => x"70",
1528 => x"3D",
1529 => x"0A",
1530 => x"6F",
1531 => x"64",
1532 => x"64",
1533 => x"00",
1534 => x"43",
1535 => x"43",
1536 => x"00",
1537 => x"07",
1538 => x"70",
1539 => x"6F",
1540 => x"64",
1541 => x"65",
1542 => x"72",
1543 => x"72",
1544 => x"3A",
1545 => x"00",
1546 => x"4F",
1547 => x"00",
1548 => x"43",
1549 => x"43",
1550 => x"42",
1551 => x"44",
1552 => x"00",
1553 => x"77",
1554 => x"74",
1555 => x"68",
1556 => x"74",
1557 => x"20",
1558 => x"65",
1559 => x"20",
1560 => x"61",
1561 => x"64",
1562 => x"72",
1563 => x"74",
1564 => x"2C",
1565 => x"74",
1566 => x"70",
1567 => x"20",
1568 => x"55",
1569 => x"20",
1570 => x"65",
1571 => x"65",
1572 => x"61",
1573 => x"20",
1574 => x"69",
1575 => x"65",
1576 => x"20",
1577 => x"6F",
1578 => x"73",
1579 => x"74",
1580 => x"20",
1581 => x"41",
1582 => x"54",
1583 => x"00",
1584 => x"65",
1585 => x"20",
1586 => x"41",
1587 => x"54",
1588 => x"73",
1589 => x"65",
1590 => x"64",
1591 => x"00",
1592 => x"45",
1593 => x"65",
1594 => x"75",
1595 => x"65",
1596 => x"00",
1597 => x"2E",
1598 => x"0A",
1599 => x"00",
1600 => x"23",
1601 => x"3A",
1602 => x"00",
1603 => x"20",
1604 => x"00",
1605 => x"08",
1606 => x"20",
1607 => x"08",
1608 => x"20",
1609 => x"20",
1610 => x"20",
1611 => x"20",
1612 => x"00",
1613 => x"00",
1614 => x"61",
1615 => x"6B",
1616 => x"77",
1617 => x"73",
1618 => x"68",
1619 => x"72",
1620 => x"2E",
1621 => x"3A",
1622 => x"29",
1623 => x"FF",
1624 => x"00",
1625 => x"00",
1626 => x"6E",
1627 => x"70",
1628 => x"20",
1629 => x"00",
1630 => x"00",
1631 => x"0F",
1632 => x"61",
1633 => x"64",
1634 => x"20",
1635 => x"00",
1636 => x"00",
1637 => x"0F",
1638 => x"61",
1639 => x"64",
1640 => x"20",
1641 => x"00",
1642 => x"00",
1643 => x"0F",
1644 => x"78",
1645 => x"72",
1646 => x"20",
1647 => x"F0",
1648 => x"00",
1649 => x"05",
1650 => x"74",
1651 => x"74",
1652 => x"6E",
1653 => x"F0",
1654 => x"40",
1655 => x"05",
1656 => x"74",
1657 => x"74",
1658 => x"7A",
1659 => x"E0",
1660 => x"80",
1661 => x"06",
1662 => x"62",
1663 => x"74",
1664 => x"6E",
1665 => x"E0",
1666 => x"C0",
1667 => x"06",
1668 => x"62",
1669 => x"74",
1670 => x"7A",
1671 => x"00",
1672 => x"00",
1673 => x"10",
1674 => x"73",
1675 => x"62",
1676 => x"6C",
1677 => x"00",
1678 => x"00",
1679 => x"0F",
1680 => x"6D",
1681 => x"6C",
1682 => x"20",
1683 => x"00",
1684 => x"00",
1685 => x"03",
1686 => x"73",
1687 => x"6D",
1688 => x"20",
1689 => x"00",
1690 => x"00",
1691 => x"0B",
1692 => x"6C",
1693 => x"62",
1694 => x"20",
1695 => x"00",
1696 => x"00",
1697 => x"04",
1698 => x"6D",
1699 => x"6D",
1700 => x"20",
1701 => x"00",
1702 => x"00",
1703 => x"0C",
1704 => x"67",
1705 => x"74",
1706 => x"63",
1707 => x"0F",
1708 => x"00",
1709 => x"07",
1710 => x"6D",
1711 => x"76",
1712 => x"20",
1713 => x"00",
1714 => x"00",
1715 => x"11",
1716 => x"69",
1717 => x"63",
1718 => x"20",
1719 => x"0F",
1720 => x"00",
1721 => x"0D",
1722 => x"6C",
1723 => x"77",
1724 => x"20",
1725 => x"0F",
1726 => x"00",
1727 => x"0E",
1728 => x"6C",
1729 => x"64",
1730 => x"20",
1731 => x"F0",
1732 => x"00",
1733 => x"01",
1734 => x"73",
1735 => x"74",
1736 => x"76",
1737 => x"FF",
1738 => x"00",
1739 => x"00",
1740 => x"72",
1741 => x"74",
1742 => x"20",
1743 => x"F0",
1744 => x"00",
1745 => x"01",
1746 => x"73",
1747 => x"74",
1748 => x"77",
1749 => x"FF",
1750 => x"00",
1751 => x"00",
1752 => x"72",
1753 => x"74",
1754 => x"20",
1755 => x"0F",
1756 => x"00",
1757 => x"02",
1758 => x"67",
1759 => x"74",
1760 => x"72",
1761 => x"0F",
1762 => x"00",
1763 => x"02",
1764 => x"67",
1765 => x"74",
1766 => x"72",
1767 => x"00",
1768 => x"00",
1769 => x"08",
1770 => x"73",
1771 => x"61",
1772 => x"62",
1773 => x"00",
1774 => x"00",
1775 => x"08",
1776 => x"73",
1777 => x"61",
1778 => x"77",
1779 => x"00",
1780 => x"00",
1781 => x"08",
1782 => x"6E",
1783 => x"74",
1784 => x"20",
1785 => x"F0",
1786 => x"00",
1787 => x"01",
1788 => x"6C",
1789 => x"6D",
1790 => x"20",
1791 => x"00",
1792 => x"00",
1793 => x"08",
1794 => x"6C",
1795 => x"72",
1796 => x"20",
1797 => x"00",
1798 => x"00",
1799 => x"08",
1800 => x"61",
1801 => x"72",
1802 => x"20",
1803 => x"F0",
1804 => x"00",
1805 => x"0A",
1806 => x"6D",
1807 => x"76",
1808 => x"20",
1809 => x"F0",
1810 => x"10",
1811 => x"0A",
1812 => x"6D",
1813 => x"76",
1814 => x"20",
1815 => x"F0",
1816 => x"20",
1817 => x"0A",
1818 => x"6D",
1819 => x"76",
1820 => x"20",
1821 => x"00",
1822 => x"00",
1823 => x"09",
1824 => x"6D",
1825 => x"76",
1826 => x"20",
1827 => x"00",
1828 => x"00",
1829 => x"09",
1830 => x"6D",
1831 => x"76",
1832 => x"20",
1833 => x"00",
1834 => x"00",
1835 => x"09",
1836 => x"6D",
1837 => x"76",
1838 => x"77",
1839 => x"00",
1840 => x"00",
1841 => x"09",
1842 => x"6D",
1843 => x"76",
1844 => x"20",
1845 => x"00",
1846 => x"00",
1847 => x"00",
1848 => x"3F",
1849 => x"3F",
1850 => x"20",
1851 => x"0F",
1852 => x"00",
1853 => x"00",
1854 => x"00",
1855 => x"00",
1856 => x"00",
1857 => x"00",
1858 => x"00",
1859 => x"00",
1860 => x"00",
1861 => x"00",
1862 => x"00",
1863 => x"00",
1864 => x"00",
1865 => x"00",
1866 => x"00",
1867 => x"00",
1868 => x"00",
1869 => x"00",
1870 => x"00",
1871 => x"00",
1872 => x"00",
1873 => x"00",
1874 => x"00",
1875 => x"00",
1876 => x"00",
1877 => x"00",
1878 => x"00",
1879 => x"00",
1880 => x"00",
1881 => x"00",
1882 => x"00",
1883 => x"00",
1884 => x"00",
1885 => x"00",
1886 => x"00",
1887 => x"00",
1888 => x"00",
1889 => x"00",
1890 => x"00",
1891 => x"00",
1892 => x"00",
1893 => x"00",
1894 => x"00",
1895 => x"00",
1896 => x"00",
1897 => x"00",
1898 => x"00",
1899 => x"00",
1900 => x"00",
1901 => x"00",
1902 => x"00",
1903 => x"00",
1904 => x"00",
1905 => x"00",
1906 => x"00",
1907 => x"00",
1908 => x"00",
1909 => x"00",
1910 => x"00",
1911 => x"00",
1912 => x"00",
1913 => x"00",
1914 => x"00",
1915 => x"00",
1916 => x"00",
1917 => x"00",
1918 => x"00",
1919 => x"00",
1920 => x"00",
1921 => x"00",
1922 => x"00",
1923 => x"00",
1924 => x"00",
1925 => x"00",
1926 => x"00",
1927 => x"00",
1928 => x"00",
1929 => x"00",
1930 => x"00",
1931 => x"00",
1932 => x"00",
1933 => x"00",
1934 => x"00",
1935 => x"00",
1936 => x"00",
1937 => x"00",
1938 => x"00",
1939 => x"00",
1940 => x"00",
1941 => x"00",
1942 => x"00",
1943 => x"00",
1944 => x"00",
1945 => x"00",
1946 => x"00",
1947 => x"00",
1948 => x"00",
1949 => x"00",
1950 => x"D1",
1951 => x"DE",


others => x"00"
);

attribute syn_ramstyle : string;
attribute syn_ramstyle of RAM : signal is "block_ram";

begin
   --busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(conv_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(conv_integer(addr_r));
end architecture behavioral; -- Entity: Sweet32_ROM